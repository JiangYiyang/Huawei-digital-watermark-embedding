`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/08/17 14:50:42
// Design Name: 
// Module Name: arctan
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module arctan(
input wire signed [40:1] y,
input wire signed [40:1] x,
output wire signed [24:1] rad

    );
wire [1:0] sig;
wire signed [40:1] y_abs;
wire signed [40:1] x_abs;
reg  signed [24:1] rad_tmp;
wire signed [40:1] y_x;
assign y_x = x == 0 ? 20000 : y_abs * 256 / x_abs; //+8
assign sig = {y[40],x[40]};
assign x_abs = x[40] ? -x : x ;
assign y_abs = y[40] ? -y : y ;
assign rad = sig[1]? ( sig[0]? (rad_tmp - 23'd6588398):(- rad_tmp)):( sig[0]? (23'd6588398-rad_tmp):(rad_tmp)) ;
always @(*) begin
 if(y_x >= 20000)
   rad_tmp =24'b001100100100001111110110;
 if(y_x > 2048 && y_x < 20000)
   rad_tmp = 15 * y_x + 40'd3000663;
 else begin

  case (y_x)
  40'd0: rad_tmp = 24'd0;
  40'd1: rad_tmp = 24'b000000000011001101111001;
  40'd2: rad_tmp = 24'b000000000110011011110010;
  40'd3: rad_tmp = 24'b000000001000000010101110;
  40'd4: rad_tmp = 24'b000000001001101001101010;
  40'd5: rad_tmp = 24'b000000001011010000100111;
  40'd6: rad_tmp = 24'b000000001110011110100000;
  40'd7: rad_tmp = 24'b000000010000000101011100;
  40'd8: rad_tmp = 24'b000000010001101100011000;
  40'd9: rad_tmp = 24'b000000010011010011010101;
  40'd10: rad_tmp = 24'b000000010110100001001110;
  40'd11: rad_tmp = 24'b000000011000001000001010;
  40'd12: rad_tmp = 24'b000000011001101111000110;
  40'd13: rad_tmp = 24'b000000011011010110000011;
  40'd14: rad_tmp = 24'b000000011110100011111100;
  40'd15: rad_tmp = 24'b000000100000001010111000;
  40'd16: rad_tmp = 24'b000000100001110001110100;
  40'd17: rad_tmp = 24'b000000100011011000110001;
  40'd18: rad_tmp = 24'b000000100100111111101101;
  40'd19: rad_tmp = 24'b000000101000001101100110;
  40'd20: rad_tmp = 24'b000000101001110100100010;
  40'd21: rad_tmp = 24'b000000101011011011011111;
  40'd22: rad_tmp = 24'b000000101101000010011011;
  40'd23: rad_tmp = 24'b000000110000010000010100;
  40'd24: rad_tmp = 24'b000000110001110111010000;
  40'd25: rad_tmp = 24'b000000110011011110001101;
  40'd26: rad_tmp = 24'b000000110101000101001001;
  40'd27: rad_tmp = 24'b000000111000010011000010;
  40'd28: rad_tmp = 24'b000000111001111001111110;
  40'd29: rad_tmp = 24'b000000111011100000111011;
  40'd30: rad_tmp = 24'b000000111101000111110111;
  40'd31: rad_tmp = 24'b000000111110101110110011;
  40'd32: rad_tmp = 24'b000001000001111100101100;
  40'd33: rad_tmp = 24'b000001000011100011101001;
  40'd34: rad_tmp = 24'b000001000101001010100101;
  40'd35: rad_tmp = 24'b000001000110110001100001;
  40'd36: rad_tmp = 24'b000001001001111111011010;
  40'd37: rad_tmp = 24'b000001001011100110010111;
  40'd38: rad_tmp = 24'b000001001101001101010011;
  40'd39: rad_tmp = 24'b000001001110110100001111;
  40'd40: rad_tmp = 24'b000001010000011011001100;
  40'd41: rad_tmp = 24'b000001010011101001000101;
  40'd42: rad_tmp = 24'b000001010101010000000001;
  40'd43: rad_tmp = 24'b000001010110110110111101;
  40'd44: rad_tmp = 24'b000001011000011101111010;
  40'd45: rad_tmp = 24'b000001011010000100110110;
  40'd46: rad_tmp = 24'b000001011101010010101111;
  40'd47: rad_tmp = 24'b000001011110111001101011;
  40'd48: rad_tmp = 24'b000001100000100000101000;
  40'd49: rad_tmp = 24'b000001100010000111100100;
  40'd50: rad_tmp = 24'b000001100011101110100001;
  40'd51: rad_tmp = 24'b000001100110111100011001;
  40'd52: rad_tmp = 24'b000001101000100011010110;
  40'd53: rad_tmp = 24'b000001101010001010010010;
  40'd54: rad_tmp = 24'b000001101011110001001111;
  40'd55: rad_tmp = 24'b000001101101011000001011;
  40'd56: rad_tmp = 24'b000001110000100110000100;
  40'd57: rad_tmp = 24'b000001110010001101000000;
  40'd58: rad_tmp = 24'b000001110011110011111101;
  40'd59: rad_tmp = 24'b000001110101011010111001;
  40'd60: rad_tmp = 24'b000001110111000001110101;
  40'd61: rad_tmp = 24'b000001111010001111101110;
  40'd62: rad_tmp = 24'b000001111011110110101011;
  40'd63: rad_tmp = 24'b000001111101011101100111;
  40'd64: rad_tmp = 24'b000001111111000100100011;
  40'd65: rad_tmp = 24'b000010000000101011100000;
  40'd66: rad_tmp = 24'b000010000010010010011100;
  40'd67: rad_tmp = 24'b000010000101100000010101;
  40'd68: rad_tmp = 24'b000010000111000111010001;
  40'd69: rad_tmp = 24'b000010001000101110001110;
  40'd70: rad_tmp = 24'b000010001010010101001010;
  40'd71: rad_tmp = 24'b000010001011111100000111;
  40'd72: rad_tmp = 24'b000010001101100011000011;
  40'd73: rad_tmp = 24'b000010001111001001111111;
  40'd74: rad_tmp = 24'b000010010010010111111000;
  40'd75: rad_tmp = 24'b000010010011111110110101;
  40'd76: rad_tmp = 24'b000010010101100101110001;
  40'd77: rad_tmp = 24'b000010010111001100101101;
  40'd78: rad_tmp = 24'b000010011000110011101010;
  40'd79: rad_tmp = 24'b000010011010011010100110;
  40'd80: rad_tmp = 24'b000010011100000001100011;
  40'd81: rad_tmp = 24'b000010011111001111011011;
  40'd82: rad_tmp = 24'b000010100000110110011000;
  40'd83: rad_tmp = 24'b000010100010011101010100;
  40'd84: rad_tmp = 24'b000010100100000100010001;
  40'd85: rad_tmp = 24'b000010100101101011001101;
  40'd86: rad_tmp = 24'b000010100111010010001001;
  40'd87: rad_tmp = 24'b000010101000111001000110;
  40'd88: rad_tmp = 24'b000010101010100000000010;
  40'd89: rad_tmp = 24'b000010101101101101111011;
  40'd90: rad_tmp = 24'b000010101111010100110111;
  40'd91: rad_tmp = 24'b000010110000111011110100;
  40'd92: rad_tmp = 24'b000010110010100010110000;
  40'd93: rad_tmp = 24'b000010110100001001101100;
  40'd94: rad_tmp = 24'b000010110101110000101001;
  40'd95: rad_tmp = 24'b000010110111010111100101;
  40'd96: rad_tmp = 24'b000010111000111110100010;
  40'd97: rad_tmp = 24'b000010111010100101011110;
  40'd98: rad_tmp = 24'b000010111100001100011010;
  40'd99: rad_tmp = 24'b000010111101110011010111;
  40'd100: rad_tmp = 24'b000011000001000001010000;
  40'd101: rad_tmp = 24'b000011000010101000001100;
  40'd102: rad_tmp = 24'b000011000100001111001000;
  40'd103: rad_tmp = 24'b000011000101110110000101;
  40'd104: rad_tmp = 24'b000011000111011101000001;
  40'd105: rad_tmp = 24'b000011001001000011111110;
  40'd106: rad_tmp = 24'b000011001010101010111010;
  40'd107: rad_tmp = 24'b000011001100010001110110;
  40'd108: rad_tmp = 24'b000011001101111000110011;
  40'd109: rad_tmp = 24'b000011001111011111101111;
  40'd110: rad_tmp = 24'b000011010001000110101100;
  40'd111: rad_tmp = 24'b000011010010101101101000;
  40'd112: rad_tmp = 24'b000011010100010100100100;
  40'd113: rad_tmp = 24'b000011010101111011100001;
  40'd114: rad_tmp = 24'b000011010111100010011101;
  40'd115: rad_tmp = 24'b000011011001001001011010;
  40'd116: rad_tmp = 24'b000011011010110000010110;
  40'd117: rad_tmp = 24'b000011011100010111010010;
  40'd118: rad_tmp = 24'b000011011101111110001111;
  40'd119: rad_tmp = 24'b000011100001001100001000;
  40'd120: rad_tmp = 24'b000011100010110011000100;
  40'd121: rad_tmp = 24'b000011100100011010000000;
  40'd122: rad_tmp = 24'b000011100110000000111101;
  40'd123: rad_tmp = 24'b000011100111100111111001;
  40'd124: rad_tmp = 24'b000011101001001110110110;
  40'd125: rad_tmp = 24'b000011101010110101110010;
  40'd126: rad_tmp = 24'b000011101100011100101110;
  40'd127: rad_tmp = 24'b000011101110000011101011;
  40'd128: rad_tmp = 24'b000011101111101010100111;
  40'd129: rad_tmp = 24'b000011110001010001100100;
  40'd130: rad_tmp = 24'b000011110010111000100000;
  40'd131: rad_tmp = 24'b000011110100011111011100;
  40'd132: rad_tmp = 24'b000011110110000110011001;
  40'd133: rad_tmp = 24'b000011110111101101010101;
  40'd134: rad_tmp = 24'b000011110111101101010101;
  40'd135: rad_tmp = 24'b000011111001010100010010;
  40'd136: rad_tmp = 24'b000011111010111011001110;
  40'd137: rad_tmp = 24'b000011111100100010001010;
  40'd138: rad_tmp = 24'b000011111110001001000111;
  40'd139: rad_tmp = 24'b000011111111110000000011;
  40'd140: rad_tmp = 24'b000100000001010111000000;
  40'd141: rad_tmp = 24'b000100000010111101111100;
  40'd142: rad_tmp = 24'b000100000100100100111000;
  40'd143: rad_tmp = 24'b000100000110001011110101;
  40'd144: rad_tmp = 24'b000100000111110010110001;
  40'd145: rad_tmp = 24'b000100001001011001101110;
  40'd146: rad_tmp = 24'b000100001011000000101010;
  40'd147: rad_tmp = 24'b000100001100100111100110;
  40'd148: rad_tmp = 24'b000100001110001110100011;
  40'd149: rad_tmp = 24'b000100001111110101011111;
  40'd150: rad_tmp = 24'b000100010001011100011100;
  40'd151: rad_tmp = 24'b000100010011000011011000;
  40'd152: rad_tmp = 24'b000100010100101010010100;
  40'd153: rad_tmp = 24'b000100010100101010010100;
  40'd154: rad_tmp = 24'b000100010110010001010001;
  40'd155: rad_tmp = 24'b000100010111111000001101;
  40'd156: rad_tmp = 24'b000100011001011111001010;
  40'd157: rad_tmp = 24'b000100011011000110000110;
  40'd158: rad_tmp = 24'b000100011100101101000010;
  40'd159: rad_tmp = 24'b000100011110010011111111;
  40'd160: rad_tmp = 24'b000100011111111010111011;
  40'd161: rad_tmp = 24'b000100100001100001111000;
  40'd162: rad_tmp = 24'b000100100011001000110100;
  40'd163: rad_tmp = 24'b000100100011001000110100;
  40'd164: rad_tmp = 24'b000100100100101111110000;
  40'd165: rad_tmp = 24'b000100100110010110101101;
  40'd166: rad_tmp = 24'b000100100111111101101001;
  40'd167: rad_tmp = 24'b000100101001100100100110;
  40'd168: rad_tmp = 24'b000100101011001011100010;
  40'd169: rad_tmp = 24'b000100101100110010011110;
  40'd170: rad_tmp = 24'b000100101110011001011011;
  40'd171: rad_tmp = 24'b000100101110011001011011;
  40'd172: rad_tmp = 24'b000100110000000000010111;
  40'd173: rad_tmp = 24'b000100110001100111010011;
  40'd174: rad_tmp = 24'b000100110011001110010000;
  40'd175: rad_tmp = 24'b000100110100110101001100;
  40'd176: rad_tmp = 24'b000100110110011100001001;
  40'd177: rad_tmp = 24'b000100110110011100001001;
  40'd178: rad_tmp = 24'b000100111000000011000101;
  40'd179: rad_tmp = 24'b000100111001101010000001;
  40'd180: rad_tmp = 24'b000100111011010000111110;
  40'd181: rad_tmp = 24'b000100111100110111111010;
  40'd182: rad_tmp = 24'b000100111110011110110111;
  40'd183: rad_tmp = 24'b000100111110011110110111;
  40'd184: rad_tmp = 24'b000101000000000101110011;
  40'd185: rad_tmp = 24'b000101000001101100101111;
  40'd186: rad_tmp = 24'b000101000011010011101100;
  40'd187: rad_tmp = 24'b000101000100111010101000;
  40'd188: rad_tmp = 24'b000101000110100001100101;
  40'd189: rad_tmp = 24'b000101000110100001100101;
  40'd190: rad_tmp = 24'b000101001000001000100001;
  40'd191: rad_tmp = 24'b000101001001101111011101;
  40'd192: rad_tmp = 24'b000101001011010110011010;
  40'd193: rad_tmp = 24'b000101001100111101010110;
  40'd194: rad_tmp = 24'b000101001100111101010110;
  40'd195: rad_tmp = 24'b000101001110100100010011;
  40'd196: rad_tmp = 24'b000101010000001011001111;
  40'd197: rad_tmp = 24'b000101010001110010001011;
  40'd198: rad_tmp = 24'b000101010001110010001011;
  40'd199: rad_tmp = 24'b000101010011011001001000;
  40'd200: rad_tmp = 24'b000101010101000000000100;
  40'd201: rad_tmp = 24'b000101010110100111000001;
  40'd202: rad_tmp = 24'b000101011000001101111101;
  40'd203: rad_tmp = 24'b000101011000001101111101;
  40'd204: rad_tmp = 24'b000101011001110100111001;
  40'd205: rad_tmp = 24'b000101011011011011110110;
  40'd206: rad_tmp = 24'b000101011101000010110010;
  40'd207: rad_tmp = 24'b000101011101000010110010;
  40'd208: rad_tmp = 24'b000101011110101001101111;
  40'd209: rad_tmp = 24'b000101100000010000101011;
  40'd210: rad_tmp = 24'b000101100001110111100111;
  40'd211: rad_tmp = 24'b000101100001110111100111;
  40'd212: rad_tmp = 24'b000101100011011110100100;
  40'd213: rad_tmp = 24'b000101100101000101100000;
  40'd214: rad_tmp = 24'b000101100101000101100000;
  40'd215: rad_tmp = 24'b000101100110101100011101;
  40'd216: rad_tmp = 24'b000101101000010011011001;
  40'd217: rad_tmp = 24'b000101101001111010010101;
  40'd218: rad_tmp = 24'b000101101001111010010101;
  40'd219: rad_tmp = 24'b000101101011100001010010;
  40'd220: rad_tmp = 24'b000101101101001000001110;
  40'd221: rad_tmp = 24'b000101101110101111001011;
  40'd222: rad_tmp = 24'b000101101110101111001011;
  40'd223: rad_tmp = 24'b000101110000010110000111;
  40'd224: rad_tmp = 24'b000101110001111101000011;
  40'd225: rad_tmp = 24'b000101110001111101000011;
  40'd226: rad_tmp = 24'b000101110011100100000000;
  40'd227: rad_tmp = 24'b000101110101001010111100;
  40'd228: rad_tmp = 24'b000101110101001010111100;
  40'd229: rad_tmp = 24'b000101110110110001111001;
  40'd230: rad_tmp = 24'b000101111000011000110101;
  40'd231: rad_tmp = 24'b000101111001111111110001;
  40'd232: rad_tmp = 24'b000101111001111111110001;
  40'd233: rad_tmp = 24'b000101111011100110101110;
  40'd234: rad_tmp = 24'b000101111101001101101010;
  40'd235: rad_tmp = 24'b000101111101001101101010;
  40'd236: rad_tmp = 24'b000101111110110100100111;
  40'd237: rad_tmp = 24'b000110000000011011100011;
  40'd238: rad_tmp = 24'b000110000000011011100011;
  40'd239: rad_tmp = 24'b000110000010000010011111;
  40'd240: rad_tmp = 24'b000110000011101001011100;
  40'd241: rad_tmp = 24'b000110000011101001011100;
  40'd242: rad_tmp = 24'b000110000101010000011000;
  40'd243: rad_tmp = 24'b000110000110110111010101;
  40'd244: rad_tmp = 24'b000110000110110111010101;
  40'd245: rad_tmp = 24'b000110001000011110010001;
  40'd246: rad_tmp = 24'b000110001000011110010001;
  40'd247: rad_tmp = 24'b000110001010000101001101;
  40'd248: rad_tmp = 24'b000110001011101100001010;
  40'd249: rad_tmp = 24'b000110001011101100001010;
  40'd250: rad_tmp = 24'b000110001101010011000110;
  40'd251: rad_tmp = 24'b000110001110111010000011;
  40'd252: rad_tmp = 24'b000110001110111010000011;
  40'd253: rad_tmp = 24'b000110010000100000111111;
  40'd254: rad_tmp = 24'b000110010010000111111011;
  40'd255: rad_tmp = 24'b000110010010000111111011;
  40'd256: rad_tmp = 24'b000110010011101110111000;
  40'd257: rad_tmp = 24'b000110010011101110111000;
  40'd258: rad_tmp = 24'b000110010101010101110100;
  40'd259: rad_tmp = 24'b000110010110111100110001;
  40'd260: rad_tmp = 24'b000110010110111100110001;
  40'd261: rad_tmp = 24'b000110011000100011101101;
  40'd262: rad_tmp = 24'b000110011000100011101101;
  40'd263: rad_tmp = 24'b000110011010001010101001;
  40'd264: rad_tmp = 24'b000110011011110001100110;
  40'd265: rad_tmp = 24'b000110011011110001100110;
  40'd266: rad_tmp = 24'b000110011101011000100010;
  40'd267: rad_tmp = 24'b000110011101011000100010;
  40'd268: rad_tmp = 24'b000110011110111111011111;
  40'd269: rad_tmp = 24'b000110100000100110011011;
  40'd270: rad_tmp = 24'b000110100000100110011011;
  40'd271: rad_tmp = 24'b000110100010001101010111;
  40'd272: rad_tmp = 24'b000110100010001101010111;
  40'd273: rad_tmp = 24'b000110100011110100010100;
  40'd274: rad_tmp = 24'b000110100101011011010000;
  40'd275: rad_tmp = 24'b000110100101011011010000;
  40'd276: rad_tmp = 24'b000110100111000010001100;
  40'd277: rad_tmp = 24'b000110100111000010001100;
  40'd278: rad_tmp = 24'b000110101000101001001001;
  40'd279: rad_tmp = 24'b000110101000101001001001;
  40'd280: rad_tmp = 24'b000110101010010000000101;
  40'd281: rad_tmp = 24'b000110101011110111000010;
  40'd282: rad_tmp = 24'b000110101011110111000010;
  40'd283: rad_tmp = 24'b000110101101011101111110;
  40'd284: rad_tmp = 24'b000110101101011101111110;
  40'd285: rad_tmp = 24'b000110101111000100111010;
  40'd286: rad_tmp = 24'b000110101111000100111010;
  40'd287: rad_tmp = 24'b000110110000101011110111;
  40'd288: rad_tmp = 24'b000110110000101011110111;
  40'd289: rad_tmp = 24'b000110110010010010110011;
  40'd290: rad_tmp = 24'b000110110011111001110000;
  40'd291: rad_tmp = 24'b000110110011111001110000;
  40'd292: rad_tmp = 24'b000110110101100000101100;
  40'd293: rad_tmp = 24'b000110110101100000101100;
  40'd294: rad_tmp = 24'b000110110111000111101000;
  40'd295: rad_tmp = 24'b000110110111000111101000;
  40'd296: rad_tmp = 24'b000110111000101110100101;
  40'd297: rad_tmp = 24'b000110111000101110100101;
  40'd298: rad_tmp = 24'b000110111010010101100001;
  40'd299: rad_tmp = 24'b000110111010010101100001;
  40'd300: rad_tmp = 24'b000110111011111100011110;
  40'd301: rad_tmp = 24'b000110111011111100011110;
  40'd302: rad_tmp = 24'b000110111101100011011010;
  40'd303: rad_tmp = 24'b000110111101100011011010;
  40'd304: rad_tmp = 24'b000110111111001010010110;
  40'd305: rad_tmp = 24'b000110111111001010010110;
  40'd306: rad_tmp = 24'b000111000000110001010011;
  40'd307: rad_tmp = 24'b000111000010011000001111;
  40'd308: rad_tmp = 24'b000111000010011000001111;
  40'd309: rad_tmp = 24'b000111000011111111001100;
  40'd310: rad_tmp = 24'b000111000011111111001100;
  40'd311: rad_tmp = 24'b000111000101100110001000;
  40'd312: rad_tmp = 24'b000111000101100110001000;
  40'd313: rad_tmp = 24'b000111000111001101000100;
  40'd314: rad_tmp = 24'b000111000111001101000100;
  40'd315: rad_tmp = 24'b000111001000110100000001;
  40'd316: rad_tmp = 24'b000111001000110100000001;
  40'd317: rad_tmp = 24'b000111001010011010111101;
  40'd318: rad_tmp = 24'b000111001010011010111101;
  40'd319: rad_tmp = 24'b000111001010011010111101;
  40'd320: rad_tmp = 24'b000111001100000001111010;
  40'd321: rad_tmp = 24'b000111001100000001111010;
  40'd322: rad_tmp = 24'b000111001101101000110110;
  40'd323: rad_tmp = 24'b000111001101101000110110;
  40'd324: rad_tmp = 24'b000111001111001111110010;
  40'd325: rad_tmp = 24'b000111001111001111110010;
  40'd326: rad_tmp = 24'b000111010000110110101111;
  40'd327: rad_tmp = 24'b000111010000110110101111;
  40'd328: rad_tmp = 24'b000111010010011101101011;
  40'd329: rad_tmp = 24'b000111010010011101101011;
  40'd330: rad_tmp = 24'b000111010100000100101000;
  40'd331: rad_tmp = 24'b000111010100000100101000;
  40'd332: rad_tmp = 24'b000111010101101011100100;
  40'd333: rad_tmp = 24'b000111010101101011100100;
  40'd334: rad_tmp = 24'b000111010111010010100000;
  40'd335: rad_tmp = 24'b000111010111010010100000;
  40'd336: rad_tmp = 24'b000111010111010010100000;
  40'd337: rad_tmp = 24'b000111011000111001011101;
  40'd338: rad_tmp = 24'b000111011000111001011101;
  40'd339: rad_tmp = 24'b000111011010100000011001;
  40'd340: rad_tmp = 24'b000111011010100000011001;
  40'd341: rad_tmp = 24'b000111011100000111010110;
  40'd342: rad_tmp = 24'b000111011100000111010110;
  40'd343: rad_tmp = 24'b000111011101101110010010;
  40'd344: rad_tmp = 24'b000111011101101110010010;
  40'd345: rad_tmp = 24'b000111011111010101001110;
  40'd346: rad_tmp = 24'b000111011111010101001110;
  40'd347: rad_tmp = 24'b000111011111010101001110;
  40'd348: rad_tmp = 24'b000111100000111100001011;
  40'd349: rad_tmp = 24'b000111100000111100001011;
  40'd350: rad_tmp = 24'b000111100010100011000111;
  40'd351: rad_tmp = 24'b000111100010100011000111;
  40'd352: rad_tmp = 24'b000111100100001010000100;
  40'd353: rad_tmp = 24'b000111100100001010000100;
  40'd354: rad_tmp = 24'b000111100100001010000100;
  40'd355: rad_tmp = 24'b000111100101110001000000;
  40'd356: rad_tmp = 24'b000111100101110001000000;
  40'd357: rad_tmp = 24'b000111100111010111111100;
  40'd358: rad_tmp = 24'b000111100111010111111100;
  40'd359: rad_tmp = 24'b000111101000111110111001;
  40'd360: rad_tmp = 24'b000111101000111110111001;
  40'd361: rad_tmp = 24'b000111101000111110111001;
  40'd362: rad_tmp = 24'b000111101010100101110101;
  40'd363: rad_tmp = 24'b000111101010100101110101;
  40'd364: rad_tmp = 24'b000111101100001100110010;
  40'd365: rad_tmp = 24'b000111101100001100110010;
  40'd366: rad_tmp = 24'b000111101100001100110010;
  40'd367: rad_tmp = 24'b000111101101110011101110;
  40'd368: rad_tmp = 24'b000111101101110011101110;
  40'd369: rad_tmp = 24'b000111101111011010101010;
  40'd370: rad_tmp = 24'b000111101111011010101010;
  40'd371: rad_tmp = 24'b000111101111011010101010;
  40'd372: rad_tmp = 24'b000111110001000001100111;
  40'd373: rad_tmp = 24'b000111110001000001100111;
  40'd374: rad_tmp = 24'b000111110010101000100011;
  40'd375: rad_tmp = 24'b000111110010101000100011;
  40'd376: rad_tmp = 24'b000111110010101000100011;
  40'd377: rad_tmp = 24'b000111110100001111100000;
  40'd378: rad_tmp = 24'b000111110100001111100000;
  40'd379: rad_tmp = 24'b000111110101110110011100;
  40'd380: rad_tmp = 24'b000111110101110110011100;
  40'd381: rad_tmp = 24'b000111110101110110011100;
  40'd382: rad_tmp = 24'b000111110111011101011000;
  40'd383: rad_tmp = 24'b000111110111011101011000;
  40'd384: rad_tmp = 24'b000111111001000100010101;
  40'd385: rad_tmp = 24'b000111111001000100010101;
  40'd386: rad_tmp = 24'b000111111001000100010101;
  40'd387: rad_tmp = 24'b000111111010101011010001;
  40'd388: rad_tmp = 24'b000111111010101011010001;
  40'd389: rad_tmp = 24'b000111111010101011010001;
  40'd390: rad_tmp = 24'b000111111100010010001110;
  40'd391: rad_tmp = 24'b000111111100010010001110;
  40'd392: rad_tmp = 24'b000111111101111001001010;
  40'd393: rad_tmp = 24'b000111111101111001001010;
  40'd394: rad_tmp = 24'b000111111101111001001010;
  40'd395: rad_tmp = 24'b000111111111100000000110;
  40'd396: rad_tmp = 24'b000111111111100000000110;
  40'd397: rad_tmp = 24'b000111111111100000000110;
  40'd398: rad_tmp = 24'b001000000001000111000011;
  40'd399: rad_tmp = 24'b001000000001000111000011;
  40'd400: rad_tmp = 24'b001000000001000111000011;
  40'd401: rad_tmp = 24'b001000000010101101111111;
  40'd402: rad_tmp = 24'b001000000010101101111111;
  40'd403: rad_tmp = 24'b001000000100010100111100;
  40'd404: rad_tmp = 24'b001000000100010100111100;
  40'd405: rad_tmp = 24'b001000000100010100111100;
  40'd406: rad_tmp = 24'b001000000101111011111000;
  40'd407: rad_tmp = 24'b001000000101111011111000;
  40'd408: rad_tmp = 24'b001000000101111011111000;
  40'd409: rad_tmp = 24'b001000000111100010110100;
  40'd410: rad_tmp = 24'b001000000111100010110100;
  40'd411: rad_tmp = 24'b001000000111100010110100;
  40'd412: rad_tmp = 24'b001000001001001001110001;
  40'd413: rad_tmp = 24'b001000001001001001110001;
  40'd414: rad_tmp = 24'b001000001001001001110001;
  40'd415: rad_tmp = 24'b001000001010110000101101;
  40'd416: rad_tmp = 24'b001000001010110000101101;
  40'd417: rad_tmp = 24'b001000001010110000101101;
  40'd418: rad_tmp = 24'b001000001100010111101010;
  40'd419: rad_tmp = 24'b001000001100010111101010;
  40'd420: rad_tmp = 24'b001000001100010111101010;
  40'd421: rad_tmp = 24'b001000001101111110100110;
  40'd422: rad_tmp = 24'b001000001101111110100110;
  40'd423: rad_tmp = 24'b001000001101111110100110;
  40'd424: rad_tmp = 24'b001000001111100101100010;
  40'd425: rad_tmp = 24'b001000001111100101100010;
  40'd426: rad_tmp = 24'b001000001111100101100010;
  40'd427: rad_tmp = 24'b001000010001001100011111;
  40'd428: rad_tmp = 24'b001000010001001100011111;
  40'd429: rad_tmp = 24'b001000010001001100011111;
  40'd430: rad_tmp = 24'b001000010010110011011011;
  40'd431: rad_tmp = 24'b001000010010110011011011;
  40'd432: rad_tmp = 24'b001000010010110011011011;
  40'd433: rad_tmp = 24'b001000010100011010011000;
  40'd434: rad_tmp = 24'b001000010100011010011000;
  40'd435: rad_tmp = 24'b001000010100011010011000;
  40'd436: rad_tmp = 24'b001000010110000001010100;
  40'd437: rad_tmp = 24'b001000010110000001010100;
  40'd438: rad_tmp = 24'b001000010110000001010100;
  40'd439: rad_tmp = 24'b001000010111101000010000;
  40'd440: rad_tmp = 24'b001000010111101000010000;
  40'd441: rad_tmp = 24'b001000010111101000010000;
  40'd442: rad_tmp = 24'b001000011001001111001101;
  40'd443: rad_tmp = 24'b001000011001001111001101;
  40'd444: rad_tmp = 24'b001000011001001111001101;
  40'd445: rad_tmp = 24'b001000011001001111001101;
  40'd446: rad_tmp = 24'b001000011010110110001001;
  40'd447: rad_tmp = 24'b001000011010110110001001;
  40'd448: rad_tmp = 24'b001000011010110110001001;
  40'd449: rad_tmp = 24'b001000011100011101000101;
  40'd450: rad_tmp = 24'b001000011100011101000101;
  40'd451: rad_tmp = 24'b001000011100011101000101;
  40'd452: rad_tmp = 24'b001000011110000100000010;
  40'd453: rad_tmp = 24'b001000011110000100000010;
  40'd454: rad_tmp = 24'b001000011110000100000010;
  40'd455: rad_tmp = 24'b001000011111101010111110;
  40'd456: rad_tmp = 24'b001000011111101010111110;
  40'd457: rad_tmp = 24'b001000011111101010111110;
  40'd458: rad_tmp = 24'b001000011111101010111110;
  40'd459: rad_tmp = 24'b001000100001010001111011;
  40'd460: rad_tmp = 24'b001000100001010001111011;
  40'd461: rad_tmp = 24'b001000100001010001111011;
  40'd462: rad_tmp = 24'b001000100010111000110111;
  40'd463: rad_tmp = 24'b001000100010111000110111;
  40'd464: rad_tmp = 24'b001000100010111000110111;
  40'd465: rad_tmp = 24'b001000100010111000110111;
  40'd466: rad_tmp = 24'b001000100100011111110011;
  40'd467: rad_tmp = 24'b001000100100011111110011;
  40'd468: rad_tmp = 24'b001000100100011111110011;
  40'd469: rad_tmp = 24'b001000100110000110110000;
  40'd470: rad_tmp = 24'b001000100110000110110000;
  40'd471: rad_tmp = 24'b001000100110000110110000;
  40'd472: rad_tmp = 24'b001000100110000110110000;
  40'd473: rad_tmp = 24'b001000100111101101101100;
  40'd474: rad_tmp = 24'b001000100111101101101100;
  40'd475: rad_tmp = 24'b001000100111101101101100;
  40'd476: rad_tmp = 24'b001000101001010100101001;
  40'd477: rad_tmp = 24'b001000101001010100101001;
  40'd478: rad_tmp = 24'b001000101001010100101001;
  40'd479: rad_tmp = 24'b001000101001010100101001;
  40'd480: rad_tmp = 24'b001000101010111011100101;
  40'd481: rad_tmp = 24'b001000101010111011100101;
  40'd482: rad_tmp = 24'b001000101010111011100101;
  40'd483: rad_tmp = 24'b001000101100100010100001;
  40'd484: rad_tmp = 24'b001000101100100010100001;
  40'd485: rad_tmp = 24'b001000101100100010100001;
  40'd486: rad_tmp = 24'b001000101100100010100001;
  40'd487: rad_tmp = 24'b001000101110001001011110;
  40'd488: rad_tmp = 24'b001000101110001001011110;
  40'd489: rad_tmp = 24'b001000101110001001011110;
  40'd490: rad_tmp = 24'b001000101110001001011110;
  40'd491: rad_tmp = 24'b001000101111110000011010;
  40'd492: rad_tmp = 24'b001000101111110000011010;
  40'd493: rad_tmp = 24'b001000101111110000011010;
  40'd494: rad_tmp = 24'b001000101111110000011010;
  40'd495: rad_tmp = 24'b001000110001010111010111;
  40'd496: rad_tmp = 24'b001000110001010111010111;
  40'd497: rad_tmp = 24'b001000110001010111010111;
  40'd498: rad_tmp = 24'b001000110001010111010111;
  40'd499: rad_tmp = 24'b001000110010111110010011;
  40'd500: rad_tmp = 24'b001000110010111110010011;
  40'd501: rad_tmp = 24'b001000110010111110010011;
  40'd502: rad_tmp = 24'b001000110100100101001111;
  40'd503: rad_tmp = 24'b001000110100100101001111;
  40'd504: rad_tmp = 24'b001000110100100101001111;
  40'd505: rad_tmp = 24'b001000110100100101001111;
  40'd506: rad_tmp = 24'b001000110110001100001100;
  40'd507: rad_tmp = 24'b001000110110001100001100;
  40'd508: rad_tmp = 24'b001000110110001100001100;
  40'd509: rad_tmp = 24'b001000110110001100001100;
  40'd510: rad_tmp = 24'b001000110111110011001000;
  40'd511: rad_tmp = 24'b001000110111110011001000;
  40'd512: rad_tmp = 24'b001000110111110011001000;
  40'd513: rad_tmp = 24'b001000110111110011001000;
  40'd514: rad_tmp = 24'b001000111001011010000101;
  40'd515: rad_tmp = 24'b001000111001011010000101;
  40'd516: rad_tmp = 24'b001000111001011010000101;
  40'd517: rad_tmp = 24'b001000111001011010000101;
  40'd518: rad_tmp = 24'b001000111011000001000001;
  40'd519: rad_tmp = 24'b001000111011000001000001;
  40'd520: rad_tmp = 24'b001000111011000001000001;
  40'd521: rad_tmp = 24'b001000111011000001000001;
  40'd522: rad_tmp = 24'b001000111011000001000001;
  40'd523: rad_tmp = 24'b001000111100100111111101;
  40'd524: rad_tmp = 24'b001000111100100111111101;
  40'd525: rad_tmp = 24'b001000111100100111111101;
  40'd526: rad_tmp = 24'b001000111100100111111101;
  40'd527: rad_tmp = 24'b001000111110001110111010;
  40'd528: rad_tmp = 24'b001000111110001110111010;
  40'd529: rad_tmp = 24'b001000111110001110111010;
  40'd530: rad_tmp = 24'b001000111110001110111010;
  40'd531: rad_tmp = 24'b001000111111110101110110;
  40'd532: rad_tmp = 24'b001000111111110101110110;
  40'd533: rad_tmp = 24'b001000111111110101110110;
  40'd534: rad_tmp = 24'b001000111111110101110110;
  40'd535: rad_tmp = 24'b001001000001011100110011;
  40'd536: rad_tmp = 24'b001001000001011100110011;
  40'd537: rad_tmp = 24'b001001000001011100110011;
  40'd538: rad_tmp = 24'b001001000001011100110011;
  40'd539: rad_tmp = 24'b001001000001011100110011;
  40'd540: rad_tmp = 24'b001001000011000011101111;
  40'd541: rad_tmp = 24'b001001000011000011101111;
  40'd542: rad_tmp = 24'b001001000011000011101111;
  40'd543: rad_tmp = 24'b001001000011000011101111;
  40'd544: rad_tmp = 24'b001001000100101010101011;
  40'd545: rad_tmp = 24'b001001000100101010101011;
  40'd546: rad_tmp = 24'b001001000100101010101011;
  40'd547: rad_tmp = 24'b001001000100101010101011;
  40'd548: rad_tmp = 24'b001001000110010001101000;
  40'd549: rad_tmp = 24'b001001000110010001101000;
  40'd550: rad_tmp = 24'b001001000110010001101000;
  40'd551: rad_tmp = 24'b001001000110010001101000;
  40'd552: rad_tmp = 24'b001001000110010001101000;
  40'd553: rad_tmp = 24'b001001000111111000100100;
  40'd554: rad_tmp = 24'b001001000111111000100100;
  40'd555: rad_tmp = 24'b001001000111111000100100;
  40'd556: rad_tmp = 24'b001001000111111000100100;
  40'd557: rad_tmp = 24'b001001000111111000100100;
  40'd558: rad_tmp = 24'b001001001001011111100001;
  40'd559: rad_tmp = 24'b001001001001011111100001;
  40'd560: rad_tmp = 24'b001001001001011111100001;
  40'd561: rad_tmp = 24'b001001001001011111100001;
  40'd562: rad_tmp = 24'b001001001011000110011101;
  40'd563: rad_tmp = 24'b001001001011000110011101;
  40'd564: rad_tmp = 24'b001001001011000110011101;
  40'd565: rad_tmp = 24'b001001001011000110011101;
  40'd566: rad_tmp = 24'b001001001011000110011101;
  40'd567: rad_tmp = 24'b001001001100101101011001;
  40'd568: rad_tmp = 24'b001001001100101101011001;
  40'd569: rad_tmp = 24'b001001001100101101011001;
  40'd570: rad_tmp = 24'b001001001100101101011001;
  40'd571: rad_tmp = 24'b001001001100101101011001;
  40'd572: rad_tmp = 24'b001001001110010100010110;
  40'd573: rad_tmp = 24'b001001001110010100010110;
  40'd574: rad_tmp = 24'b001001001110010100010110;
  40'd575: rad_tmp = 24'b001001001110010100010110;
  40'd576: rad_tmp = 24'b001001001110010100010110;
  40'd577: rad_tmp = 24'b001001001111111011010010;
  40'd578: rad_tmp = 24'b001001001111111011010010;
  40'd579: rad_tmp = 24'b001001001111111011010010;
  40'd580: rad_tmp = 24'b001001001111111011010010;
  40'd581: rad_tmp = 24'b001001001111111011010010;
  40'd582: rad_tmp = 24'b001001010001100010001111;
  40'd583: rad_tmp = 24'b001001010001100010001111;
  40'd584: rad_tmp = 24'b001001010001100010001111;
  40'd585: rad_tmp = 24'b001001010001100010001111;
  40'd586: rad_tmp = 24'b001001010001100010001111;
  40'd587: rad_tmp = 24'b001001010011001001001011;
  40'd588: rad_tmp = 24'b001001010011001001001011;
  40'd589: rad_tmp = 24'b001001010011001001001011;
  40'd590: rad_tmp = 24'b001001010011001001001011;
  40'd591: rad_tmp = 24'b001001010011001001001011;
  40'd592: rad_tmp = 24'b001001010100110000000111;
  40'd593: rad_tmp = 24'b001001010100110000000111;
  40'd594: rad_tmp = 24'b001001010100110000000111;
  40'd595: rad_tmp = 24'b001001010100110000000111;
  40'd596: rad_tmp = 24'b001001010100110000000111;
  40'd597: rad_tmp = 24'b001001010110010111000100;
  40'd598: rad_tmp = 24'b001001010110010111000100;
  40'd599: rad_tmp = 24'b001001010110010111000100;
  40'd600: rad_tmp = 24'b001001010110010111000100;
  40'd601: rad_tmp = 24'b001001010110010111000100;
  40'd602: rad_tmp = 24'b001001010111111110000000;
  40'd603: rad_tmp = 24'b001001010111111110000000;
  40'd604: rad_tmp = 24'b001001010111111110000000;
  40'd605: rad_tmp = 24'b001001010111111110000000;
  40'd606: rad_tmp = 24'b001001010111111110000000;
  40'd607: rad_tmp = 24'b001001011001100100111101;
  40'd608: rad_tmp = 24'b001001011001100100111101;
  40'd609: rad_tmp = 24'b001001011001100100111101;
  40'd610: rad_tmp = 24'b001001011001100100111101;
  40'd611: rad_tmp = 24'b001001011001100100111101;
  40'd612: rad_tmp = 24'b001001011001100100111101;
  40'd613: rad_tmp = 24'b001001011011001011111001;
  40'd614: rad_tmp = 24'b001001011011001011111001;
  40'd615: rad_tmp = 24'b001001011011001011111001;
  40'd616: rad_tmp = 24'b001001011011001011111001;
  40'd617: rad_tmp = 24'b001001011011001011111001;
  40'd618: rad_tmp = 24'b001001011100110010110101;
  40'd619: rad_tmp = 24'b001001011100110010110101;
  40'd620: rad_tmp = 24'b001001011100110010110101;
  40'd621: rad_tmp = 24'b001001011100110010110101;
  40'd622: rad_tmp = 24'b001001011100110010110101;
  40'd623: rad_tmp = 24'b001001011100110010110101;
  40'd624: rad_tmp = 24'b001001011110011001110010;
  40'd625: rad_tmp = 24'b001001011110011001110010;
  40'd626: rad_tmp = 24'b001001011110011001110010;
  40'd627: rad_tmp = 24'b001001011110011001110010;
  40'd628: rad_tmp = 24'b001001011110011001110010;
  40'd629: rad_tmp = 24'b001001100000000000101110;
  40'd630: rad_tmp = 24'b001001100000000000101110;
  40'd631: rad_tmp = 24'b001001100000000000101110;
  40'd632: rad_tmp = 24'b001001100000000000101110;
  40'd633: rad_tmp = 24'b001001100000000000101110;
  40'd634: rad_tmp = 24'b001001100000000000101110;
  40'd635: rad_tmp = 24'b001001100001100111101011;
  40'd636: rad_tmp = 24'b001001100001100111101011;
  40'd637: rad_tmp = 24'b001001100001100111101011;
  40'd638: rad_tmp = 24'b001001100001100111101011;
  40'd639: rad_tmp = 24'b001001100001100111101011;
  40'd640: rad_tmp = 24'b001001100001100111101011;
  40'd641: rad_tmp = 24'b001001100011001110100111;
  40'd642: rad_tmp = 24'b001001100011001110100111;
  40'd643: rad_tmp = 24'b001001100011001110100111;
  40'd644: rad_tmp = 24'b001001100011001110100111;
  40'd645: rad_tmp = 24'b001001100011001110100111;
  40'd646: rad_tmp = 24'b001001100011001110100111;
  40'd647: rad_tmp = 24'b001001100100110101100011;
  40'd648: rad_tmp = 24'b001001100100110101100011;
  40'd649: rad_tmp = 24'b001001100100110101100011;
  40'd650: rad_tmp = 24'b001001100100110101100011;
  40'd651: rad_tmp = 24'b001001100100110101100011;
  40'd652: rad_tmp = 24'b001001100100110101100011;
  40'd653: rad_tmp = 24'b001001100110011100100000;
  40'd654: rad_tmp = 24'b001001100110011100100000;
  40'd655: rad_tmp = 24'b001001100110011100100000;
  40'd656: rad_tmp = 24'b001001100110011100100000;
  40'd657: rad_tmp = 24'b001001100110011100100000;
  40'd658: rad_tmp = 24'b001001100110011100100000;
  40'd659: rad_tmp = 24'b001001101000000011011100;
  40'd660: rad_tmp = 24'b001001101000000011011100;
  40'd661: rad_tmp = 24'b001001101000000011011100;
  40'd662: rad_tmp = 24'b001001101000000011011100;
  40'd663: rad_tmp = 24'b001001101000000011011100;
  40'd664: rad_tmp = 24'b001001101000000011011100;
  40'd665: rad_tmp = 24'b001001101001101010011001;
  40'd666: rad_tmp = 24'b001001101001101010011001;
  40'd667: rad_tmp = 24'b001001101001101010011001;
  40'd668: rad_tmp = 24'b001001101001101010011001;
  40'd669: rad_tmp = 24'b001001101001101010011001;
  40'd670: rad_tmp = 24'b001001101001101010011001;
  40'd671: rad_tmp = 24'b001001101011010001010101;
  40'd672: rad_tmp = 24'b001001101011010001010101;
  40'd673: rad_tmp = 24'b001001101011010001010101;
  40'd674: rad_tmp = 24'b001001101011010001010101;
  40'd675: rad_tmp = 24'b001001101011010001010101;
  40'd676: rad_tmp = 24'b001001101011010001010101;
  40'd677: rad_tmp = 24'b001001101100111000010001;
  40'd678: rad_tmp = 24'b001001101100111000010001;
  40'd679: rad_tmp = 24'b001001101100111000010001;
  40'd680: rad_tmp = 24'b001001101100111000010001;
  40'd681: rad_tmp = 24'b001001101100111000010001;
  40'd682: rad_tmp = 24'b001001101100111000010001;
  40'd683: rad_tmp = 24'b001001101100111000010001;
  40'd684: rad_tmp = 24'b001001101110011111001110;
  40'd685: rad_tmp = 24'b001001101110011111001110;
  40'd686: rad_tmp = 24'b001001101110011111001110;
  40'd687: rad_tmp = 24'b001001101110011111001110;
  40'd688: rad_tmp = 24'b001001101110011111001110;
  40'd689: rad_tmp = 24'b001001101110011111001110;
  40'd690: rad_tmp = 24'b001001101110011111001110;
  40'd691: rad_tmp = 24'b001001110000000110001010;
  40'd692: rad_tmp = 24'b001001110000000110001010;
  40'd693: rad_tmp = 24'b001001110000000110001010;
  40'd694: rad_tmp = 24'b001001110000000110001010;
  40'd695: rad_tmp = 24'b001001110000000110001010;
  40'd696: rad_tmp = 24'b001001110000000110001010;
  40'd697: rad_tmp = 24'b001001110001101101000111;
  40'd698: rad_tmp = 24'b001001110001101101000111;
  40'd699: rad_tmp = 24'b001001110001101101000111;
  40'd700: rad_tmp = 24'b001001110001101101000111;
  40'd701: rad_tmp = 24'b001001110001101101000111;
  40'd702: rad_tmp = 24'b001001110001101101000111;
  40'd703: rad_tmp = 24'b001001110001101101000111;
  40'd704: rad_tmp = 24'b001001110011010100000011;
  40'd705: rad_tmp = 24'b001001110011010100000011;
  40'd706: rad_tmp = 24'b001001110011010100000011;
  40'd707: rad_tmp = 24'b001001110011010100000011;
  40'd708: rad_tmp = 24'b001001110011010100000011;
  40'd709: rad_tmp = 24'b001001110011010100000011;
  40'd710: rad_tmp = 24'b001001110011010100000011;
  40'd711: rad_tmp = 24'b001001110100111010111111;
  40'd712: rad_tmp = 24'b001001110100111010111111;
  40'd713: rad_tmp = 24'b001001110100111010111111;
  40'd714: rad_tmp = 24'b001001110100111010111111;
  40'd715: rad_tmp = 24'b001001110100111010111111;
  40'd716: rad_tmp = 24'b001001110100111010111111;
  40'd717: rad_tmp = 24'b001001110100111010111111;
  40'd718: rad_tmp = 24'b001001110110100001111100;
  40'd719: rad_tmp = 24'b001001110110100001111100;
  40'd720: rad_tmp = 24'b001001110110100001111100;
  40'd721: rad_tmp = 24'b001001110110100001111100;
  40'd722: rad_tmp = 24'b001001110110100001111100;
  40'd723: rad_tmp = 24'b001001110110100001111100;
  40'd724: rad_tmp = 24'b001001110110100001111100;
  40'd725: rad_tmp = 24'b001001111000001000111000;
  40'd726: rad_tmp = 24'b001001111000001000111000;
  40'd727: rad_tmp = 24'b001001111000001000111000;
  40'd728: rad_tmp = 24'b001001111000001000111000;
  40'd729: rad_tmp = 24'b001001111000001000111000;
  40'd730: rad_tmp = 24'b001001111000001000111000;
  40'd731: rad_tmp = 24'b001001111000001000111000;
  40'd732: rad_tmp = 24'b001001111000001000111000;
  40'd733: rad_tmp = 24'b001001111001101111110101;
  40'd734: rad_tmp = 24'b001001111001101111110101;
  40'd735: rad_tmp = 24'b001001111001101111110101;
  40'd736: rad_tmp = 24'b001001111001101111110101;
  40'd737: rad_tmp = 24'b001001111001101111110101;
  40'd738: rad_tmp = 24'b001001111001101111110101;
  40'd739: rad_tmp = 24'b001001111001101111110101;
  40'd740: rad_tmp = 24'b001001111011010110110001;
  40'd741: rad_tmp = 24'b001001111011010110110001;
  40'd742: rad_tmp = 24'b001001111011010110110001;
  40'd743: rad_tmp = 24'b001001111011010110110001;
  40'd744: rad_tmp = 24'b001001111011010110110001;
  40'd745: rad_tmp = 24'b001001111011010110110001;
  40'd746: rad_tmp = 24'b001001111011010110110001;
  40'd747: rad_tmp = 24'b001001111011010110110001;
  40'd748: rad_tmp = 24'b001001111100111101101101;
  40'd749: rad_tmp = 24'b001001111100111101101101;
  40'd750: rad_tmp = 24'b001001111100111101101101;
  40'd751: rad_tmp = 24'b001001111100111101101101;
  40'd752: rad_tmp = 24'b001001111100111101101101;
  40'd753: rad_tmp = 24'b001001111100111101101101;
  40'd754: rad_tmp = 24'b001001111100111101101101;
  40'd755: rad_tmp = 24'b001001111110100100101010;
  40'd756: rad_tmp = 24'b001001111110100100101010;
  40'd757: rad_tmp = 24'b001001111110100100101010;
  40'd758: rad_tmp = 24'b001001111110100100101010;
  40'd759: rad_tmp = 24'b001001111110100100101010;
  40'd760: rad_tmp = 24'b001001111110100100101010;
  40'd761: rad_tmp = 24'b001001111110100100101010;
  40'd762: rad_tmp = 24'b001001111110100100101010;
  40'd763: rad_tmp = 24'b001010000000001011100110;
  40'd764: rad_tmp = 24'b001010000000001011100110;
  40'd765: rad_tmp = 24'b001010000000001011100110;
  40'd766: rad_tmp = 24'b001010000000001011100110;
  40'd767: rad_tmp = 24'b001010000000001011100110;
  40'd768: rad_tmp = 24'b001010000000001011100110;
  40'd769: rad_tmp = 24'b001010000000001011100110;
  40'd770: rad_tmp = 24'b001010000000001011100110;
  40'd771: rad_tmp = 24'b001010000001110010100011;
  40'd772: rad_tmp = 24'b001010000001110010100011;
  40'd773: rad_tmp = 24'b001010000001110010100011;
  40'd774: rad_tmp = 24'b001010000001110010100011;
  40'd775: rad_tmp = 24'b001010000001110010100011;
  40'd776: rad_tmp = 24'b001010000001110010100011;
  40'd777: rad_tmp = 24'b001010000001110010100011;
  40'd778: rad_tmp = 24'b001010000001110010100011;
  40'd779: rad_tmp = 24'b001010000001110010100011;
  40'd780: rad_tmp = 24'b001010000011011001011111;
  40'd781: rad_tmp = 24'b001010000011011001011111;
  40'd782: rad_tmp = 24'b001010000011011001011111;
  40'd783: rad_tmp = 24'b001010000011011001011111;
  40'd784: rad_tmp = 24'b001010000011011001011111;
  40'd785: rad_tmp = 24'b001010000011011001011111;
  40'd786: rad_tmp = 24'b001010000011011001011111;
  40'd787: rad_tmp = 24'b001010000011011001011111;
  40'd788: rad_tmp = 24'b001010000101000000011011;
  40'd789: rad_tmp = 24'b001010000101000000011011;
  40'd790: rad_tmp = 24'b001010000101000000011011;
  40'd791: rad_tmp = 24'b001010000101000000011011;
  40'd792: rad_tmp = 24'b001010000101000000011011;
  40'd793: rad_tmp = 24'b001010000101000000011011;
  40'd794: rad_tmp = 24'b001010000101000000011011;
  40'd795: rad_tmp = 24'b001010000101000000011011;
  40'd796: rad_tmp = 24'b001010000110100111011000;
  40'd797: rad_tmp = 24'b001010000110100111011000;
  40'd798: rad_tmp = 24'b001010000110100111011000;
  40'd799: rad_tmp = 24'b001010000110100111011000;
  40'd800: rad_tmp = 24'b001010000110100111011000;
  40'd801: rad_tmp = 24'b001010000110100111011000;
  40'd802: rad_tmp = 24'b001010000110100111011000;
  40'd803: rad_tmp = 24'b001010000110100111011000;
  40'd804: rad_tmp = 24'b001010000110100111011000;
  40'd805: rad_tmp = 24'b001010001000001110010100;
  40'd806: rad_tmp = 24'b001010001000001110010100;
  40'd807: rad_tmp = 24'b001010001000001110010100;
  40'd808: rad_tmp = 24'b001010001000001110010100;
  40'd809: rad_tmp = 24'b001010001000001110010100;
  40'd810: rad_tmp = 24'b001010001000001110010100;
  40'd811: rad_tmp = 24'b001010001000001110010100;
  40'd812: rad_tmp = 24'b001010001000001110010100;
  40'd813: rad_tmp = 24'b001010001000001110010100;
  40'd814: rad_tmp = 24'b001010001001110101010001;
  40'd815: rad_tmp = 24'b001010001001110101010001;
  40'd816: rad_tmp = 24'b001010001001110101010001;
  40'd817: rad_tmp = 24'b001010001001110101010001;
  40'd818: rad_tmp = 24'b001010001001110101010001;
  40'd819: rad_tmp = 24'b001010001001110101010001;
  40'd820: rad_tmp = 24'b001010001001110101010001;
  40'd821: rad_tmp = 24'b001010001001110101010001;
  40'd822: rad_tmp = 24'b001010001001110101010001;
  40'd823: rad_tmp = 24'b001010001011011100001101;
  40'd824: rad_tmp = 24'b001010001011011100001101;
  40'd825: rad_tmp = 24'b001010001011011100001101;
  40'd826: rad_tmp = 24'b001010001011011100001101;
  40'd827: rad_tmp = 24'b001010001011011100001101;
  40'd828: rad_tmp = 24'b001010001011011100001101;
  40'd829: rad_tmp = 24'b001010001011011100001101;
  40'd830: rad_tmp = 24'b001010001011011100001101;
  40'd831: rad_tmp = 24'b001010001011011100001101;
  40'd832: rad_tmp = 24'b001010001101000011001001;
  40'd833: rad_tmp = 24'b001010001101000011001001;
  40'd834: rad_tmp = 24'b001010001101000011001001;
  40'd835: rad_tmp = 24'b001010001101000011001001;
  40'd836: rad_tmp = 24'b001010001101000011001001;
  40'd837: rad_tmp = 24'b001010001101000011001001;
  40'd838: rad_tmp = 24'b001010001101000011001001;
  40'd839: rad_tmp = 24'b001010001101000011001001;
  40'd840: rad_tmp = 24'b001010001101000011001001;
  40'd841: rad_tmp = 24'b001010001101000011001001;
  40'd842: rad_tmp = 24'b001010001110101010000110;
  40'd843: rad_tmp = 24'b001010001110101010000110;
  40'd844: rad_tmp = 24'b001010001110101010000110;
  40'd845: rad_tmp = 24'b001010001110101010000110;
  40'd846: rad_tmp = 24'b001010001110101010000110;
  40'd847: rad_tmp = 24'b001010001110101010000110;
  40'd848: rad_tmp = 24'b001010001110101010000110;
  40'd849: rad_tmp = 24'b001010001110101010000110;
  40'd850: rad_tmp = 24'b001010001110101010000110;
  40'd851: rad_tmp = 24'b001010010000010001000010;
  40'd852: rad_tmp = 24'b001010010000010001000010;
  40'd853: rad_tmp = 24'b001010010000010001000010;
  40'd854: rad_tmp = 24'b001010010000010001000010;
  40'd855: rad_tmp = 24'b001010010000010001000010;
  40'd856: rad_tmp = 24'b001010010000010001000010;
  40'd857: rad_tmp = 24'b001010010000010001000010;
  40'd858: rad_tmp = 24'b001010010000010001000010;
  40'd859: rad_tmp = 24'b001010010000010001000010;
  40'd860: rad_tmp = 24'b001010010000010001000010;
  40'd861: rad_tmp = 24'b001010010001110111111111;
  40'd862: rad_tmp = 24'b001010010001110111111111;
  40'd863: rad_tmp = 24'b001010010001110111111111;
  40'd864: rad_tmp = 24'b001010010001110111111111;
  40'd865: rad_tmp = 24'b001010010001110111111111;
  40'd866: rad_tmp = 24'b001010010001110111111111;
  40'd867: rad_tmp = 24'b001010010001110111111111;
  40'd868: rad_tmp = 24'b001010010001110111111111;
  40'd869: rad_tmp = 24'b001010010001110111111111;
  40'd870: rad_tmp = 24'b001010010001110111111111;
  40'd871: rad_tmp = 24'b001010010011011110111011;
  40'd872: rad_tmp = 24'b001010010011011110111011;
  40'd873: rad_tmp = 24'b001010010011011110111011;
  40'd874: rad_tmp = 24'b001010010011011110111011;
  40'd875: rad_tmp = 24'b001010010011011110111011;
  40'd876: rad_tmp = 24'b001010010011011110111011;
  40'd877: rad_tmp = 24'b001010010011011110111011;
  40'd878: rad_tmp = 24'b001010010011011110111011;
  40'd879: rad_tmp = 24'b001010010011011110111011;
  40'd880: rad_tmp = 24'b001010010011011110111011;
  40'd881: rad_tmp = 24'b001010010101000101110111;
  40'd882: rad_tmp = 24'b001010010101000101110111;
  40'd883: rad_tmp = 24'b001010010101000101110111;
  40'd884: rad_tmp = 24'b001010010101000101110111;
  40'd885: rad_tmp = 24'b001010010101000101110111;
  40'd886: rad_tmp = 24'b001010010101000101110111;
  40'd887: rad_tmp = 24'b001010010101000101110111;
  40'd888: rad_tmp = 24'b001010010101000101110111;
  40'd889: rad_tmp = 24'b001010010101000101110111;
  40'd890: rad_tmp = 24'b001010010101000101110111;
  40'd891: rad_tmp = 24'b001010010101000101110111;
  40'd892: rad_tmp = 24'b001010010110101100110100;
  40'd893: rad_tmp = 24'b001010010110101100110100;
  40'd894: rad_tmp = 24'b001010010110101100110100;
  40'd895: rad_tmp = 24'b001010010110101100110100;
  40'd896: rad_tmp = 24'b001010010110101100110100;
  40'd897: rad_tmp = 24'b001010010110101100110100;
  40'd898: rad_tmp = 24'b001010010110101100110100;
  40'd899: rad_tmp = 24'b001010010110101100110100;
  40'd900: rad_tmp = 24'b001010010110101100110100;
  40'd901: rad_tmp = 24'b001010010110101100110100;
  40'd902: rad_tmp = 24'b001010011000010011110000;
  40'd903: rad_tmp = 24'b001010011000010011110000;
  40'd904: rad_tmp = 24'b001010011000010011110000;
  40'd905: rad_tmp = 24'b001010011000010011110000;
  40'd906: rad_tmp = 24'b001010011000010011110000;
  40'd907: rad_tmp = 24'b001010011000010011110000;
  40'd908: rad_tmp = 24'b001010011000010011110000;
  40'd909: rad_tmp = 24'b001010011000010011110000;
  40'd910: rad_tmp = 24'b001010011000010011110000;
  40'd911: rad_tmp = 24'b001010011000010011110000;
  40'd912: rad_tmp = 24'b001010011000010011110000;
  40'd913: rad_tmp = 24'b001010011001111010101100;
  40'd914: rad_tmp = 24'b001010011001111010101100;
  40'd915: rad_tmp = 24'b001010011001111010101100;
  40'd916: rad_tmp = 24'b001010011001111010101100;
  40'd917: rad_tmp = 24'b001010011001111010101100;
  40'd918: rad_tmp = 24'b001010011001111010101100;
  40'd919: rad_tmp = 24'b001010011001111010101100;
  40'd920: rad_tmp = 24'b001010011001111010101100;
  40'd921: rad_tmp = 24'b001010011001111010101100;
  40'd922: rad_tmp = 24'b001010011001111010101100;
  40'd923: rad_tmp = 24'b001010011001111010101100;
  40'd924: rad_tmp = 24'b001010011011100001101001;
  40'd925: rad_tmp = 24'b001010011011100001101001;
  40'd926: rad_tmp = 24'b001010011011100001101001;
  40'd927: rad_tmp = 24'b001010011011100001101001;
  40'd928: rad_tmp = 24'b001010011011100001101001;
  40'd929: rad_tmp = 24'b001010011011100001101001;
  40'd930: rad_tmp = 24'b001010011011100001101001;
  40'd931: rad_tmp = 24'b001010011011100001101001;
  40'd932: rad_tmp = 24'b001010011011100001101001;
  40'd933: rad_tmp = 24'b001010011011100001101001;
  40'd934: rad_tmp = 24'b001010011011100001101001;
  40'd935: rad_tmp = 24'b001010011011100001101001;
  40'd936: rad_tmp = 24'b001010011101001000100101;
  40'd937: rad_tmp = 24'b001010011101001000100101;
  40'd938: rad_tmp = 24'b001010011101001000100101;
  40'd939: rad_tmp = 24'b001010011101001000100101;
  40'd940: rad_tmp = 24'b001010011101001000100101;
  40'd941: rad_tmp = 24'b001010011101001000100101;
  40'd942: rad_tmp = 24'b001010011101001000100101;
  40'd943: rad_tmp = 24'b001010011101001000100101;
  40'd944: rad_tmp = 24'b001010011101001000100101;
  40'd945: rad_tmp = 24'b001010011101001000100101;
  40'd946: rad_tmp = 24'b001010011101001000100101;
  40'd947: rad_tmp = 24'b001010011110101111100010;
  40'd948: rad_tmp = 24'b001010011110101111100010;
  40'd949: rad_tmp = 24'b001010011110101111100010;
  40'd950: rad_tmp = 24'b001010011110101111100010;
  40'd951: rad_tmp = 24'b001010011110101111100010;
  40'd952: rad_tmp = 24'b001010011110101111100010;
  40'd953: rad_tmp = 24'b001010011110101111100010;
  40'd954: rad_tmp = 24'b001010011110101111100010;
  40'd955: rad_tmp = 24'b001010011110101111100010;
  40'd956: rad_tmp = 24'b001010011110101111100010;
  40'd957: rad_tmp = 24'b001010011110101111100010;
  40'd958: rad_tmp = 24'b001010011110101111100010;
  40'd959: rad_tmp = 24'b001010100000010110011110;
  40'd960: rad_tmp = 24'b001010100000010110011110;
  40'd961: rad_tmp = 24'b001010100000010110011110;
  40'd962: rad_tmp = 24'b001010100000010110011110;
  40'd963: rad_tmp = 24'b001010100000010110011110;
  40'd964: rad_tmp = 24'b001010100000010110011110;
  40'd965: rad_tmp = 24'b001010100000010110011110;
  40'd966: rad_tmp = 24'b001010100000010110011110;
  40'd967: rad_tmp = 24'b001010100000010110011110;
  40'd968: rad_tmp = 24'b001010100000010110011110;
  40'd969: rad_tmp = 24'b001010100000010110011110;
  40'd970: rad_tmp = 24'b001010100000010110011110;
  40'd971: rad_tmp = 24'b001010100000010110011110;
  40'd972: rad_tmp = 24'b001010100001111101011010;
  40'd973: rad_tmp = 24'b001010100001111101011010;
  40'd974: rad_tmp = 24'b001010100001111101011010;
  40'd975: rad_tmp = 24'b001010100001111101011010;
  40'd976: rad_tmp = 24'b001010100001111101011010;
  40'd977: rad_tmp = 24'b001010100001111101011010;
  40'd978: rad_tmp = 24'b001010100001111101011010;
  40'd979: rad_tmp = 24'b001010100001111101011010;
  40'd980: rad_tmp = 24'b001010100001111101011010;
  40'd981: rad_tmp = 24'b001010100001111101011010;
  40'd982: rad_tmp = 24'b001010100001111101011010;
  40'd983: rad_tmp = 24'b001010100001111101011010;
  40'd984: rad_tmp = 24'b001010100011100100010111;
  40'd985: rad_tmp = 24'b001010100011100100010111;
  40'd986: rad_tmp = 24'b001010100011100100010111;
  40'd987: rad_tmp = 24'b001010100011100100010111;
  40'd988: rad_tmp = 24'b001010100011100100010111;
  40'd989: rad_tmp = 24'b001010100011100100010111;
  40'd990: rad_tmp = 24'b001010100011100100010111;
  40'd991: rad_tmp = 24'b001010100011100100010111;
  40'd992: rad_tmp = 24'b001010100011100100010111;
  40'd993: rad_tmp = 24'b001010100011100100010111;
  40'd994: rad_tmp = 24'b001010100011100100010111;
  40'd995: rad_tmp = 24'b001010100011100100010111;
  40'd996: rad_tmp = 24'b001010100011100100010111;
  40'd997: rad_tmp = 24'b001010100101001011010011;
  40'd998: rad_tmp = 24'b001010100101001011010011;
  40'd999: rad_tmp = 24'b001010100101001011010011;
  40'd1000: rad_tmp = 24'b001010100101001011010011;
  40'd1001: rad_tmp = 24'b001010100101001011010011;
  40'd1002: rad_tmp = 24'b001010100101001011010011;
  40'd1003: rad_tmp = 24'b001010100101001011010011;
  40'd1004: rad_tmp = 24'b001010100101001011010011;
  40'd1005: rad_tmp = 24'b001010100101001011010011;
  40'd1006: rad_tmp = 24'b001010100101001011010011;
  40'd1007: rad_tmp = 24'b001010100101001011010011;
  40'd1008: rad_tmp = 24'b001010100101001011010011;
  40'd1009: rad_tmp = 24'b001010100101001011010011;
  40'd1010: rad_tmp = 24'b001010100110110010010000;
  40'd1011: rad_tmp = 24'b001010100110110010010000;
  40'd1012: rad_tmp = 24'b001010100110110010010000;
  40'd1013: rad_tmp = 24'b001010100110110010010000;
  40'd1014: rad_tmp = 24'b001010100110110010010000;
  40'd1015: rad_tmp = 24'b001010100110110010010000;
  40'd1016: rad_tmp = 24'b001010100110110010010000;
  40'd1017: rad_tmp = 24'b001010100110110010010000;
  40'd1018: rad_tmp = 24'b001010100110110010010000;
  40'd1019: rad_tmp = 24'b001010100110110010010000;
  40'd1020: rad_tmp = 24'b001010100110110010010000;
  40'd1021: rad_tmp = 24'b001010100110110010010000;
  40'd1022: rad_tmp = 24'b001010100110110010010000;
  40'd1023: rad_tmp = 24'b001010100110110010010000;
  40'd1024: rad_tmp = 24'b001010101000011001001100;
  40'd1025: rad_tmp = 24'b001010101000011001001100;
  40'd1026: rad_tmp = 24'b001010101000011001001100;
  40'd1027: rad_tmp = 24'b001010101000011001001100;
  40'd1028: rad_tmp = 24'b001010101000011001001100;
  40'd1029: rad_tmp = 24'b001010101000011001001100;
  40'd1030: rad_tmp = 24'b001010101000011001001100;
  40'd1031: rad_tmp = 24'b001010101000011001001100;
  40'd1032: rad_tmp = 24'b001010101000011001001100;
  40'd1033: rad_tmp = 24'b001010101000011001001100;
  40'd1034: rad_tmp = 24'b001010101000011001001100;
  40'd1035: rad_tmp = 24'b001010101000011001001100;
  40'd1036: rad_tmp = 24'b001010101000011001001100;
  40'd1037: rad_tmp = 24'b001010101000011001001100;
  40'd1038: rad_tmp = 24'b001010101010000000001000;
  40'd1039: rad_tmp = 24'b001010101010000000001000;
  40'd1040: rad_tmp = 24'b001010101010000000001000;
  40'd1041: rad_tmp = 24'b001010101010000000001000;
  40'd1042: rad_tmp = 24'b001010101010000000001000;
  40'd1043: rad_tmp = 24'b001010101010000000001000;
  40'd1044: rad_tmp = 24'b001010101010000000001000;
  40'd1045: rad_tmp = 24'b001010101010000000001000;
  40'd1046: rad_tmp = 24'b001010101010000000001000;
  40'd1047: rad_tmp = 24'b001010101010000000001000;
  40'd1048: rad_tmp = 24'b001010101010000000001000;
  40'd1049: rad_tmp = 24'b001010101010000000001000;
  40'd1050: rad_tmp = 24'b001010101010000000001000;
  40'd1051: rad_tmp = 24'b001010101010000000001000;
  40'd1052: rad_tmp = 24'b001010101011100111000101;
  40'd1053: rad_tmp = 24'b001010101011100111000101;
  40'd1054: rad_tmp = 24'b001010101011100111000101;
  40'd1055: rad_tmp = 24'b001010101011100111000101;
  40'd1056: rad_tmp = 24'b001010101011100111000101;
  40'd1057: rad_tmp = 24'b001010101011100111000101;
  40'd1058: rad_tmp = 24'b001010101011100111000101;
  40'd1059: rad_tmp = 24'b001010101011100111000101;
  40'd1060: rad_tmp = 24'b001010101011100111000101;
  40'd1061: rad_tmp = 24'b001010101011100111000101;
  40'd1062: rad_tmp = 24'b001010101011100111000101;
  40'd1063: rad_tmp = 24'b001010101011100111000101;
  40'd1064: rad_tmp = 24'b001010101011100111000101;
  40'd1065: rad_tmp = 24'b001010101011100111000101;
  40'd1066: rad_tmp = 24'b001010101101001110000001;
  40'd1067: rad_tmp = 24'b001010101101001110000001;
  40'd1068: rad_tmp = 24'b001010101101001110000001;
  40'd1069: rad_tmp = 24'b001010101101001110000001;
  40'd1070: rad_tmp = 24'b001010101101001110000001;
  40'd1071: rad_tmp = 24'b001010101101001110000001;
  40'd1072: rad_tmp = 24'b001010101101001110000001;
  40'd1073: rad_tmp = 24'b001010101101001110000001;
  40'd1074: rad_tmp = 24'b001010101101001110000001;
  40'd1075: rad_tmp = 24'b001010101101001110000001;
  40'd1076: rad_tmp = 24'b001010101101001110000001;
  40'd1077: rad_tmp = 24'b001010101101001110000001;
  40'd1078: rad_tmp = 24'b001010101101001110000001;
  40'd1079: rad_tmp = 24'b001010101101001110000001;
  40'd1080: rad_tmp = 24'b001010101101001110000001;
  40'd1081: rad_tmp = 24'b001010101110110100111110;
  40'd1082: rad_tmp = 24'b001010101110110100111110;
  40'd1083: rad_tmp = 24'b001010101110110100111110;
  40'd1084: rad_tmp = 24'b001010101110110100111110;
  40'd1085: rad_tmp = 24'b001010101110110100111110;
  40'd1086: rad_tmp = 24'b001010101110110100111110;
  40'd1087: rad_tmp = 24'b001010101110110100111110;
  40'd1088: rad_tmp = 24'b001010101110110100111110;
  40'd1089: rad_tmp = 24'b001010101110110100111110;
  40'd1090: rad_tmp = 24'b001010101110110100111110;
  40'd1091: rad_tmp = 24'b001010101110110100111110;
  40'd1092: rad_tmp = 24'b001010101110110100111110;
  40'd1093: rad_tmp = 24'b001010101110110100111110;
  40'd1094: rad_tmp = 24'b001010101110110100111110;
  40'd1095: rad_tmp = 24'b001010101110110100111110;
  40'd1096: rad_tmp = 24'b001010101110110100111110;
  40'd1097: rad_tmp = 24'b001010110000011011111010;
  40'd1098: rad_tmp = 24'b001010110000011011111010;
  40'd1099: rad_tmp = 24'b001010110000011011111010;
  40'd1100: rad_tmp = 24'b001010110000011011111010;
  40'd1101: rad_tmp = 24'b001010110000011011111010;
  40'd1102: rad_tmp = 24'b001010110000011011111010;
  40'd1103: rad_tmp = 24'b001010110000011011111010;
  40'd1104: rad_tmp = 24'b001010110000011011111010;
  40'd1105: rad_tmp = 24'b001010110000011011111010;
  40'd1106: rad_tmp = 24'b001010110000011011111010;
  40'd1107: rad_tmp = 24'b001010110000011011111010;
  40'd1108: rad_tmp = 24'b001010110000011011111010;
  40'd1109: rad_tmp = 24'b001010110000011011111010;
  40'd1110: rad_tmp = 24'b001010110000011011111010;
  40'd1111: rad_tmp = 24'b001010110000011011111010;
  40'd1112: rad_tmp = 24'b001010110010000010110110;
  40'd1113: rad_tmp = 24'b001010110010000010110110;
  40'd1114: rad_tmp = 24'b001010110010000010110110;
  40'd1115: rad_tmp = 24'b001010110010000010110110;
  40'd1116: rad_tmp = 24'b001010110010000010110110;
  40'd1117: rad_tmp = 24'b001010110010000010110110;
  40'd1118: rad_tmp = 24'b001010110010000010110110;
  40'd1119: rad_tmp = 24'b001010110010000010110110;
  40'd1120: rad_tmp = 24'b001010110010000010110110;
  40'd1121: rad_tmp = 24'b001010110010000010110110;
  40'd1122: rad_tmp = 24'b001010110010000010110110;
  40'd1123: rad_tmp = 24'b001010110010000010110110;
  40'd1124: rad_tmp = 24'b001010110010000010110110;
  40'd1125: rad_tmp = 24'b001010110010000010110110;
  40'd1126: rad_tmp = 24'b001010110010000010110110;
  40'd1127: rad_tmp = 24'b001010110010000010110110;
  40'd1128: rad_tmp = 24'b001010110010000010110110;
  40'd1129: rad_tmp = 24'b001010110011101001110011;
  40'd1130: rad_tmp = 24'b001010110011101001110011;
  40'd1131: rad_tmp = 24'b001010110011101001110011;
  40'd1132: rad_tmp = 24'b001010110011101001110011;
  40'd1133: rad_tmp = 24'b001010110011101001110011;
  40'd1134: rad_tmp = 24'b001010110011101001110011;
  40'd1135: rad_tmp = 24'b001010110011101001110011;
  40'd1136: rad_tmp = 24'b001010110011101001110011;
  40'd1137: rad_tmp = 24'b001010110011101001110011;
  40'd1138: rad_tmp = 24'b001010110011101001110011;
  40'd1139: rad_tmp = 24'b001010110011101001110011;
  40'd1140: rad_tmp = 24'b001010110011101001110011;
  40'd1141: rad_tmp = 24'b001010110011101001110011;
  40'd1142: rad_tmp = 24'b001010110011101001110011;
  40'd1143: rad_tmp = 24'b001010110011101001110011;
  40'd1144: rad_tmp = 24'b001010110011101001110011;
  40'd1145: rad_tmp = 24'b001010110101010000101111;
  40'd1146: rad_tmp = 24'b001010110101010000101111;
  40'd1147: rad_tmp = 24'b001010110101010000101111;
  40'd1148: rad_tmp = 24'b001010110101010000101111;
  40'd1149: rad_tmp = 24'b001010110101010000101111;
  40'd1150: rad_tmp = 24'b001010110101010000101111;
  40'd1151: rad_tmp = 24'b001010110101010000101111;
  40'd1152: rad_tmp = 24'b001010110101010000101111;
  40'd1153: rad_tmp = 24'b001010110101010000101111;
  40'd1154: rad_tmp = 24'b001010110101010000101111;
  40'd1155: rad_tmp = 24'b001010110101010000101111;
  40'd1156: rad_tmp = 24'b001010110101010000101111;
  40'd1157: rad_tmp = 24'b001010110101010000101111;
  40'd1158: rad_tmp = 24'b001010110101010000101111;
  40'd1159: rad_tmp = 24'b001010110101010000101111;
  40'd1160: rad_tmp = 24'b001010110101010000101111;
  40'd1161: rad_tmp = 24'b001010110101010000101111;
  40'd1162: rad_tmp = 24'b001010110110110111101100;
  40'd1163: rad_tmp = 24'b001010110110110111101100;
  40'd1164: rad_tmp = 24'b001010110110110111101100;
  40'd1165: rad_tmp = 24'b001010110110110111101100;
  40'd1166: rad_tmp = 24'b001010110110110111101100;
  40'd1167: rad_tmp = 24'b001010110110110111101100;
  40'd1168: rad_tmp = 24'b001010110110110111101100;
  40'd1169: rad_tmp = 24'b001010110110110111101100;
  40'd1170: rad_tmp = 24'b001010110110110111101100;
  40'd1171: rad_tmp = 24'b001010110110110111101100;
  40'd1172: rad_tmp = 24'b001010110110110111101100;
  40'd1173: rad_tmp = 24'b001010110110110111101100;
  40'd1174: rad_tmp = 24'b001010110110110111101100;
  40'd1175: rad_tmp = 24'b001010110110110111101100;
  40'd1176: rad_tmp = 24'b001010110110110111101100;
  40'd1177: rad_tmp = 24'b001010110110110111101100;
  40'd1178: rad_tmp = 24'b001010110110110111101100;
  40'd1179: rad_tmp = 24'b001010110110110111101100;
  40'd1180: rad_tmp = 24'b001010111000011110101000;
  40'd1181: rad_tmp = 24'b001010111000011110101000;
  40'd1182: rad_tmp = 24'b001010111000011110101000;
  40'd1183: rad_tmp = 24'b001010111000011110101000;
  40'd1184: rad_tmp = 24'b001010111000011110101000;
  40'd1185: rad_tmp = 24'b001010111000011110101000;
  40'd1186: rad_tmp = 24'b001010111000011110101000;
  40'd1187: rad_tmp = 24'b001010111000011110101000;
  40'd1188: rad_tmp = 24'b001010111000011110101000;
  40'd1189: rad_tmp = 24'b001010111000011110101000;
  40'd1190: rad_tmp = 24'b001010111000011110101000;
  40'd1191: rad_tmp = 24'b001010111000011110101000;
  40'd1192: rad_tmp = 24'b001010111000011110101000;
  40'd1193: rad_tmp = 24'b001010111000011110101000;
  40'd1194: rad_tmp = 24'b001010111000011110101000;
  40'd1195: rad_tmp = 24'b001010111000011110101000;
  40'd1196: rad_tmp = 24'b001010111000011110101000;
  40'd1197: rad_tmp = 24'b001010111000011110101000;
  40'd1198: rad_tmp = 24'b001010111010000101100100;
  40'd1199: rad_tmp = 24'b001010111010000101100100;
  40'd1200: rad_tmp = 24'b001010111010000101100100;
  40'd1201: rad_tmp = 24'b001010111010000101100100;
  40'd1202: rad_tmp = 24'b001010111010000101100100;
  40'd1203: rad_tmp = 24'b001010111010000101100100;
  40'd1204: rad_tmp = 24'b001010111010000101100100;
  40'd1205: rad_tmp = 24'b001010111010000101100100;
  40'd1206: rad_tmp = 24'b001010111010000101100100;
  40'd1207: rad_tmp = 24'b001010111010000101100100;
  40'd1208: rad_tmp = 24'b001010111010000101100100;
  40'd1209: rad_tmp = 24'b001010111010000101100100;
  40'd1210: rad_tmp = 24'b001010111010000101100100;
  40'd1211: rad_tmp = 24'b001010111010000101100100;
  40'd1212: rad_tmp = 24'b001010111010000101100100;
  40'd1213: rad_tmp = 24'b001010111010000101100100;
  40'd1214: rad_tmp = 24'b001010111010000101100100;
  40'd1215: rad_tmp = 24'b001010111010000101100100;
  40'd1216: rad_tmp = 24'b001010111010000101100100;
  40'd1217: rad_tmp = 24'b001010111011101100100001;
  40'd1218: rad_tmp = 24'b001010111011101100100001;
  40'd1219: rad_tmp = 24'b001010111011101100100001;
  40'd1220: rad_tmp = 24'b001010111011101100100001;
  40'd1221: rad_tmp = 24'b001010111011101100100001;
  40'd1222: rad_tmp = 24'b001010111011101100100001;
  40'd1223: rad_tmp = 24'b001010111011101100100001;
  40'd1224: rad_tmp = 24'b001010111011101100100001;
  40'd1225: rad_tmp = 24'b001010111011101100100001;
  40'd1226: rad_tmp = 24'b001010111011101100100001;
  40'd1227: rad_tmp = 24'b001010111011101100100001;
  40'd1228: rad_tmp = 24'b001010111011101100100001;
  40'd1229: rad_tmp = 24'b001010111011101100100001;
  40'd1230: rad_tmp = 24'b001010111011101100100001;
  40'd1231: rad_tmp = 24'b001010111011101100100001;
  40'd1232: rad_tmp = 24'b001010111011101100100001;
  40'd1233: rad_tmp = 24'b001010111011101100100001;
  40'd1234: rad_tmp = 24'b001010111011101100100001;
  40'd1235: rad_tmp = 24'b001010111011101100100001;
  40'd1236: rad_tmp = 24'b001010111101010011011101;
  40'd1237: rad_tmp = 24'b001010111101010011011101;
  40'd1238: rad_tmp = 24'b001010111101010011011101;
  40'd1239: rad_tmp = 24'b001010111101010011011101;
  40'd1240: rad_tmp = 24'b001010111101010011011101;
  40'd1241: rad_tmp = 24'b001010111101010011011101;
  40'd1242: rad_tmp = 24'b001010111101010011011101;
  40'd1243: rad_tmp = 24'b001010111101010011011101;
  40'd1244: rad_tmp = 24'b001010111101010011011101;
  40'd1245: rad_tmp = 24'b001010111101010011011101;
  40'd1246: rad_tmp = 24'b001010111101010011011101;
  40'd1247: rad_tmp = 24'b001010111101010011011101;
  40'd1248: rad_tmp = 24'b001010111101010011011101;
  40'd1249: rad_tmp = 24'b001010111101010011011101;
  40'd1250: rad_tmp = 24'b001010111101010011011101;
  40'd1251: rad_tmp = 24'b001010111101010011011101;
  40'd1252: rad_tmp = 24'b001010111101010011011101;
  40'd1253: rad_tmp = 24'b001010111101010011011101;
  40'd1254: rad_tmp = 24'b001010111101010011011101;
  40'd1255: rad_tmp = 24'b001010111101010011011101;
  40'd1256: rad_tmp = 24'b001010111110111010011010;
  40'd1257: rad_tmp = 24'b001010111110111010011010;
  40'd1258: rad_tmp = 24'b001010111110111010011010;
  40'd1259: rad_tmp = 24'b001010111110111010011010;
  40'd1260: rad_tmp = 24'b001010111110111010011010;
  40'd1261: rad_tmp = 24'b001010111110111010011010;
  40'd1262: rad_tmp = 24'b001010111110111010011010;
  40'd1263: rad_tmp = 24'b001010111110111010011010;
  40'd1264: rad_tmp = 24'b001010111110111010011010;
  40'd1265: rad_tmp = 24'b001010111110111010011010;
  40'd1266: rad_tmp = 24'b001010111110111010011010;
  40'd1267: rad_tmp = 24'b001010111110111010011010;
  40'd1268: rad_tmp = 24'b001010111110111010011010;
  40'd1269: rad_tmp = 24'b001010111110111010011010;
  40'd1270: rad_tmp = 24'b001010111110111010011010;
  40'd1271: rad_tmp = 24'b001010111110111010011010;
  40'd1272: rad_tmp = 24'b001010111110111010011010;
  40'd1273: rad_tmp = 24'b001010111110111010011010;
  40'd1274: rad_tmp = 24'b001010111110111010011010;
  40'd1275: rad_tmp = 24'b001010111110111010011010;
  40'd1276: rad_tmp = 24'b001010111110111010011010;
  40'd1277: rad_tmp = 24'b001011000000100001010110;
  40'd1278: rad_tmp = 24'b001011000000100001010110;
  40'd1279: rad_tmp = 24'b001011000000100001010110;
  40'd1280: rad_tmp = 24'b001011000000100001010110;
  40'd1281: rad_tmp = 24'b001011000000100001010110;
  40'd1282: rad_tmp = 24'b001011000000100001010110;
  40'd1283: rad_tmp = 24'b001011000000100001010110;
  40'd1284: rad_tmp = 24'b001011000000100001010110;
  40'd1285: rad_tmp = 24'b001011000000100001010110;
  40'd1286: rad_tmp = 24'b001011000000100001010110;
  40'd1287: rad_tmp = 24'b001011000000100001010110;
  40'd1288: rad_tmp = 24'b001011000000100001010110;
  40'd1289: rad_tmp = 24'b001011000000100001010110;
  40'd1290: rad_tmp = 24'b001011000000100001010110;
  40'd1291: rad_tmp = 24'b001011000000100001010110;
  40'd1292: rad_tmp = 24'b001011000000100001010110;
  40'd1293: rad_tmp = 24'b001011000000100001010110;
  40'd1294: rad_tmp = 24'b001011000000100001010110;
  40'd1295: rad_tmp = 24'b001011000000100001010110;
  40'd1296: rad_tmp = 24'b001011000000100001010110;
  40'd1297: rad_tmp = 24'b001011000000100001010110;
  40'd1298: rad_tmp = 24'b001011000010001000010010;
  40'd1299: rad_tmp = 24'b001011000010001000010010;
  40'd1300: rad_tmp = 24'b001011000010001000010010;
  40'd1301: rad_tmp = 24'b001011000010001000010010;
  40'd1302: rad_tmp = 24'b001011000010001000010010;
  40'd1303: rad_tmp = 24'b001011000010001000010010;
  40'd1304: rad_tmp = 24'b001011000010001000010010;
  40'd1305: rad_tmp = 24'b001011000010001000010010;
  40'd1306: rad_tmp = 24'b001011000010001000010010;
  40'd1307: rad_tmp = 24'b001011000010001000010010;
  40'd1308: rad_tmp = 24'b001011000010001000010010;
  40'd1309: rad_tmp = 24'b001011000010001000010010;
  40'd1310: rad_tmp = 24'b001011000010001000010010;
  40'd1311: rad_tmp = 24'b001011000010001000010010;
  40'd1312: rad_tmp = 24'b001011000010001000010010;
  40'd1313: rad_tmp = 24'b001011000010001000010010;
  40'd1314: rad_tmp = 24'b001011000010001000010010;
  40'd1315: rad_tmp = 24'b001011000010001000010010;
  40'd1316: rad_tmp = 24'b001011000010001000010010;
  40'd1317: rad_tmp = 24'b001011000010001000010010;
  40'd1318: rad_tmp = 24'b001011000010001000010010;
  40'd1319: rad_tmp = 24'b001011000011101111001111;
  40'd1320: rad_tmp = 24'b001011000011101111001111;
  40'd1321: rad_tmp = 24'b001011000011101111001111;
  40'd1322: rad_tmp = 24'b001011000011101111001111;
  40'd1323: rad_tmp = 24'b001011000011101111001111;
  40'd1324: rad_tmp = 24'b001011000011101111001111;
  40'd1325: rad_tmp = 24'b001011000011101111001111;
  40'd1326: rad_tmp = 24'b001011000011101111001111;
  40'd1327: rad_tmp = 24'b001011000011101111001111;
  40'd1328: rad_tmp = 24'b001011000011101111001111;
  40'd1329: rad_tmp = 24'b001011000011101111001111;
  40'd1330: rad_tmp = 24'b001011000011101111001111;
  40'd1331: rad_tmp = 24'b001011000011101111001111;
  40'd1332: rad_tmp = 24'b001011000011101111001111;
  40'd1333: rad_tmp = 24'b001011000011101111001111;
  40'd1334: rad_tmp = 24'b001011000011101111001111;
  40'd1335: rad_tmp = 24'b001011000011101111001111;
  40'd1336: rad_tmp = 24'b001011000011101111001111;
  40'd1337: rad_tmp = 24'b001011000011101111001111;
  40'd1338: rad_tmp = 24'b001011000011101111001111;
  40'd1339: rad_tmp = 24'b001011000011101111001111;
  40'd1340: rad_tmp = 24'b001011000011101111001111;
  40'd1341: rad_tmp = 24'b001011000011101111001111;
  40'd1342: rad_tmp = 24'b001011000101010110001011;
  40'd1343: rad_tmp = 24'b001011000101010110001011;
  40'd1344: rad_tmp = 24'b001011000101010110001011;
  40'd1345: rad_tmp = 24'b001011000101010110001011;
  40'd1346: rad_tmp = 24'b001011000101010110001011;
  40'd1347: rad_tmp = 24'b001011000101010110001011;
  40'd1348: rad_tmp = 24'b001011000101010110001011;
  40'd1349: rad_tmp = 24'b001011000101010110001011;
  40'd1350: rad_tmp = 24'b001011000101010110001011;
  40'd1351: rad_tmp = 24'b001011000101010110001011;
  40'd1352: rad_tmp = 24'b001011000101010110001011;
  40'd1353: rad_tmp = 24'b001011000101010110001011;
  40'd1354: rad_tmp = 24'b001011000101010110001011;
  40'd1355: rad_tmp = 24'b001011000101010110001011;
  40'd1356: rad_tmp = 24'b001011000101010110001011;
  40'd1357: rad_tmp = 24'b001011000101010110001011;
  40'd1358: rad_tmp = 24'b001011000101010110001011;
  40'd1359: rad_tmp = 24'b001011000101010110001011;
  40'd1360: rad_tmp = 24'b001011000101010110001011;
  40'd1361: rad_tmp = 24'b001011000101010110001011;
  40'd1362: rad_tmp = 24'b001011000101010110001011;
  40'd1363: rad_tmp = 24'b001011000101010110001011;
  40'd1364: rad_tmp = 24'b001011000101010110001011;
  40'd1365: rad_tmp = 24'b001011000110111101001000;
  40'd1366: rad_tmp = 24'b001011000110111101001000;
  40'd1367: rad_tmp = 24'b001011000110111101001000;
  40'd1368: rad_tmp = 24'b001011000110111101001000;
  40'd1369: rad_tmp = 24'b001011000110111101001000;
  40'd1370: rad_tmp = 24'b001011000110111101001000;
  40'd1371: rad_tmp = 24'b001011000110111101001000;
  40'd1372: rad_tmp = 24'b001011000110111101001000;
  40'd1373: rad_tmp = 24'b001011000110111101001000;
  40'd1374: rad_tmp = 24'b001011000110111101001000;
  40'd1375: rad_tmp = 24'b001011000110111101001000;
  40'd1376: rad_tmp = 24'b001011000110111101001000;
  40'd1377: rad_tmp = 24'b001011000110111101001000;
  40'd1378: rad_tmp = 24'b001011000110111101001000;
  40'd1379: rad_tmp = 24'b001011000110111101001000;
  40'd1380: rad_tmp = 24'b001011000110111101001000;
  40'd1381: rad_tmp = 24'b001011000110111101001000;
  40'd1382: rad_tmp = 24'b001011000110111101001000;
  40'd1383: rad_tmp = 24'b001011000110111101001000;
  40'd1384: rad_tmp = 24'b001011000110111101001000;
  40'd1385: rad_tmp = 24'b001011000110111101001000;
  40'd1386: rad_tmp = 24'b001011000110111101001000;
  40'd1387: rad_tmp = 24'b001011000110111101001000;
  40'd1388: rad_tmp = 24'b001011000110111101001000;
  40'd1389: rad_tmp = 24'b001011001000100100000100;
  40'd1390: rad_tmp = 24'b001011001000100100000100;
  40'd1391: rad_tmp = 24'b001011001000100100000100;
  40'd1392: rad_tmp = 24'b001011001000100100000100;
  40'd1393: rad_tmp = 24'b001011001000100100000100;
  40'd1394: rad_tmp = 24'b001011001000100100000100;
  40'd1395: rad_tmp = 24'b001011001000100100000100;
  40'd1396: rad_tmp = 24'b001011001000100100000100;
  40'd1397: rad_tmp = 24'b001011001000100100000100;
  40'd1398: rad_tmp = 24'b001011001000100100000100;
  40'd1399: rad_tmp = 24'b001011001000100100000100;
  40'd1400: rad_tmp = 24'b001011001000100100000100;
  40'd1401: rad_tmp = 24'b001011001000100100000100;
  40'd1402: rad_tmp = 24'b001011001000100100000100;
  40'd1403: rad_tmp = 24'b001011001000100100000100;
  40'd1404: rad_tmp = 24'b001011001000100100000100;
  40'd1405: rad_tmp = 24'b001011001000100100000100;
  40'd1406: rad_tmp = 24'b001011001000100100000100;
  40'd1407: rad_tmp = 24'b001011001000100100000100;
  40'd1408: rad_tmp = 24'b001011001000100100000100;
  40'd1409: rad_tmp = 24'b001011001000100100000100;
  40'd1410: rad_tmp = 24'b001011001000100100000100;
  40'd1411: rad_tmp = 24'b001011001000100100000100;
  40'd1412: rad_tmp = 24'b001011001000100100000100;
  40'd1413: rad_tmp = 24'b001011001000100100000100;
  40'd1414: rad_tmp = 24'b001011001010001011000000;
  40'd1415: rad_tmp = 24'b001011001010001011000000;
  40'd1416: rad_tmp = 24'b001011001010001011000000;
  40'd1417: rad_tmp = 24'b001011001010001011000000;
  40'd1418: rad_tmp = 24'b001011001010001011000000;
  40'd1419: rad_tmp = 24'b001011001010001011000000;
  40'd1420: rad_tmp = 24'b001011001010001011000000;
  40'd1421: rad_tmp = 24'b001011001010001011000000;
  40'd1422: rad_tmp = 24'b001011001010001011000000;
  40'd1423: rad_tmp = 24'b001011001010001011000000;
  40'd1424: rad_tmp = 24'b001011001010001011000000;
  40'd1425: rad_tmp = 24'b001011001010001011000000;
  40'd1426: rad_tmp = 24'b001011001010001011000000;
  40'd1427: rad_tmp = 24'b001011001010001011000000;
  40'd1428: rad_tmp = 24'b001011001010001011000000;
  40'd1429: rad_tmp = 24'b001011001010001011000000;
  40'd1430: rad_tmp = 24'b001011001010001011000000;
  40'd1431: rad_tmp = 24'b001011001010001011000000;
  40'd1432: rad_tmp = 24'b001011001010001011000000;
  40'd1433: rad_tmp = 24'b001011001010001011000000;
  40'd1434: rad_tmp = 24'b001011001010001011000000;
  40'd1435: rad_tmp = 24'b001011001010001011000000;
  40'd1436: rad_tmp = 24'b001011001010001011000000;
  40'd1437: rad_tmp = 24'b001011001010001011000000;
  40'd1438: rad_tmp = 24'b001011001010001011000000;
  40'd1439: rad_tmp = 24'b001011001010001011000000;
  40'd1440: rad_tmp = 24'b001011001011110001111101;
  40'd1441: rad_tmp = 24'b001011001011110001111101;
  40'd1442: rad_tmp = 24'b001011001011110001111101;
  40'd1443: rad_tmp = 24'b001011001011110001111101;
  40'd1444: rad_tmp = 24'b001011001011110001111101;
  40'd1445: rad_tmp = 24'b001011001011110001111101;
  40'd1446: rad_tmp = 24'b001011001011110001111101;
  40'd1447: rad_tmp = 24'b001011001011110001111101;
  40'd1448: rad_tmp = 24'b001011001011110001111101;
  40'd1449: rad_tmp = 24'b001011001011110001111101;
  40'd1450: rad_tmp = 24'b001011001011110001111101;
  40'd1451: rad_tmp = 24'b001011001011110001111101;
  40'd1452: rad_tmp = 24'b001011001011110001111101;
  40'd1453: rad_tmp = 24'b001011001011110001111101;
  40'd1454: rad_tmp = 24'b001011001011110001111101;
  40'd1455: rad_tmp = 24'b001011001011110001111101;
  40'd1456: rad_tmp = 24'b001011001011110001111101;
  40'd1457: rad_tmp = 24'b001011001011110001111101;
  40'd1458: rad_tmp = 24'b001011001011110001111101;
  40'd1459: rad_tmp = 24'b001011001011110001111101;
  40'd1460: rad_tmp = 24'b001011001011110001111101;
  40'd1461: rad_tmp = 24'b001011001011110001111101;
  40'd1462: rad_tmp = 24'b001011001011110001111101;
  40'd1463: rad_tmp = 24'b001011001011110001111101;
  40'd1464: rad_tmp = 24'b001011001011110001111101;
  40'd1465: rad_tmp = 24'b001011001011110001111101;
  40'd1466: rad_tmp = 24'b001011001011110001111101;
  40'd1467: rad_tmp = 24'b001011001101011000111001;
  40'd1468: rad_tmp = 24'b001011001101011000111001;
  40'd1469: rad_tmp = 24'b001011001101011000111001;
  40'd1470: rad_tmp = 24'b001011001101011000111001;
  40'd1471: rad_tmp = 24'b001011001101011000111001;
  40'd1472: rad_tmp = 24'b001011001101011000111001;
  40'd1473: rad_tmp = 24'b001011001101011000111001;
  40'd1474: rad_tmp = 24'b001011001101011000111001;
  40'd1475: rad_tmp = 24'b001011001101011000111001;
  40'd1476: rad_tmp = 24'b001011001101011000111001;
  40'd1477: rad_tmp = 24'b001011001101011000111001;
  40'd1478: rad_tmp = 24'b001011001101011000111001;
  40'd1479: rad_tmp = 24'b001011001101011000111001;
  40'd1480: rad_tmp = 24'b001011001101011000111001;
  40'd1481: rad_tmp = 24'b001011001101011000111001;
  40'd1482: rad_tmp = 24'b001011001101011000111001;
  40'd1483: rad_tmp = 24'b001011001101011000111001;
  40'd1484: rad_tmp = 24'b001011001101011000111001;
  40'd1485: rad_tmp = 24'b001011001101011000111001;
  40'd1486: rad_tmp = 24'b001011001101011000111001;
  40'd1487: rad_tmp = 24'b001011001101011000111001;
  40'd1488: rad_tmp = 24'b001011001101011000111001;
  40'd1489: rad_tmp = 24'b001011001101011000111001;
  40'd1490: rad_tmp = 24'b001011001101011000111001;
  40'd1491: rad_tmp = 24'b001011001101011000111001;
  40'd1492: rad_tmp = 24'b001011001101011000111001;
  40'd1493: rad_tmp = 24'b001011001101011000111001;
  40'd1494: rad_tmp = 24'b001011001101011000111001;
  40'd1495: rad_tmp = 24'b001011001110111111110110;
  40'd1496: rad_tmp = 24'b001011001110111111110110;
  40'd1497: rad_tmp = 24'b001011001110111111110110;
  40'd1498: rad_tmp = 24'b001011001110111111110110;
  40'd1499: rad_tmp = 24'b001011001110111111110110;
  40'd1500: rad_tmp = 24'b001011001110111111110110;
  40'd1501: rad_tmp = 24'b001011001110111111110110;
  40'd1502: rad_tmp = 24'b001011001110111111110110;
  40'd1503: rad_tmp = 24'b001011001110111111110110;
  40'd1504: rad_tmp = 24'b001011001110111111110110;
  40'd1505: rad_tmp = 24'b001011001110111111110110;
  40'd1506: rad_tmp = 24'b001011001110111111110110;
  40'd1507: rad_tmp = 24'b001011001110111111110110;
  40'd1508: rad_tmp = 24'b001011001110111111110110;
  40'd1509: rad_tmp = 24'b001011001110111111110110;
  40'd1510: rad_tmp = 24'b001011001110111111110110;
  40'd1511: rad_tmp = 24'b001011001110111111110110;
  40'd1512: rad_tmp = 24'b001011001110111111110110;
  40'd1513: rad_tmp = 24'b001011001110111111110110;
  40'd1514: rad_tmp = 24'b001011001110111111110110;
  40'd1515: rad_tmp = 24'b001011001110111111110110;
  40'd1516: rad_tmp = 24'b001011001110111111110110;
  40'd1517: rad_tmp = 24'b001011001110111111110110;
  40'd1518: rad_tmp = 24'b001011001110111111110110;
  40'd1519: rad_tmp = 24'b001011001110111111110110;
  40'd1520: rad_tmp = 24'b001011001110111111110110;
  40'd1521: rad_tmp = 24'b001011001110111111110110;
  40'd1522: rad_tmp = 24'b001011001110111111110110;
  40'd1523: rad_tmp = 24'b001011010000100110110010;
  40'd1524: rad_tmp = 24'b001011010000100110110010;
  40'd1525: rad_tmp = 24'b001011010000100110110010;
  40'd1526: rad_tmp = 24'b001011010000100110110010;
  40'd1527: rad_tmp = 24'b001011010000100110110010;
  40'd1528: rad_tmp = 24'b001011010000100110110010;
  40'd1529: rad_tmp = 24'b001011010000100110110010;
  40'd1530: rad_tmp = 24'b001011010000100110110010;
  40'd1531: rad_tmp = 24'b001011010000100110110010;
  40'd1532: rad_tmp = 24'b001011010000100110110010;
  40'd1533: rad_tmp = 24'b001011010000100110110010;
  40'd1534: rad_tmp = 24'b001011010000100110110010;
  40'd1535: rad_tmp = 24'b001011010000100110110010;
  40'd1536: rad_tmp = 24'b001011010000100110110010;
  40'd1537: rad_tmp = 24'b001011010000100110110010;
  40'd1538: rad_tmp = 24'b001011010000100110110010;
  40'd1539: rad_tmp = 24'b001011010000100110110010;
  40'd1540: rad_tmp = 24'b001011010000100110110010;
  40'd1541: rad_tmp = 24'b001011010000100110110010;
  40'd1542: rad_tmp = 24'b001011010000100110110010;
  40'd1543: rad_tmp = 24'b001011010000100110110010;
  40'd1544: rad_tmp = 24'b001011010000100110110010;
  40'd1545: rad_tmp = 24'b001011010000100110110010;
  40'd1546: rad_tmp = 24'b001011010000100110110010;
  40'd1547: rad_tmp = 24'b001011010000100110110010;
  40'd1548: rad_tmp = 24'b001011010000100110110010;
  40'd1549: rad_tmp = 24'b001011010000100110110010;
  40'd1550: rad_tmp = 24'b001011010000100110110010;
  40'd1551: rad_tmp = 24'b001011010000100110110010;
  40'd1552: rad_tmp = 24'b001011010000100110110010;
  40'd1553: rad_tmp = 24'b001011010010001101101110;
  40'd1554: rad_tmp = 24'b001011010010001101101110;
  40'd1555: rad_tmp = 24'b001011010010001101101110;
  40'd1556: rad_tmp = 24'b001011010010001101101110;
  40'd1557: rad_tmp = 24'b001011010010001101101110;
  40'd1558: rad_tmp = 24'b001011010010001101101110;
  40'd1559: rad_tmp = 24'b001011010010001101101110;
  40'd1560: rad_tmp = 24'b001011010010001101101110;
  40'd1561: rad_tmp = 24'b001011010010001101101110;
  40'd1562: rad_tmp = 24'b001011010010001101101110;
  40'd1563: rad_tmp = 24'b001011010010001101101110;
  40'd1564: rad_tmp = 24'b001011010010001101101110;
  40'd1565: rad_tmp = 24'b001011010010001101101110;
  40'd1566: rad_tmp = 24'b001011010010001101101110;
  40'd1567: rad_tmp = 24'b001011010010001101101110;
  40'd1568: rad_tmp = 24'b001011010010001101101110;
  40'd1569: rad_tmp = 24'b001011010010001101101110;
  40'd1570: rad_tmp = 24'b001011010010001101101110;
  40'd1571: rad_tmp = 24'b001011010010001101101110;
  40'd1572: rad_tmp = 24'b001011010010001101101110;
  40'd1573: rad_tmp = 24'b001011010010001101101110;
  40'd1574: rad_tmp = 24'b001011010010001101101110;
  40'd1575: rad_tmp = 24'b001011010010001101101110;
  40'd1576: rad_tmp = 24'b001011010010001101101110;
  40'd1577: rad_tmp = 24'b001011010010001101101110;
  40'd1578: rad_tmp = 24'b001011010010001101101110;
  40'd1579: rad_tmp = 24'b001011010010001101101110;
  40'd1580: rad_tmp = 24'b001011010010001101101110;
  40'd1581: rad_tmp = 24'b001011010010001101101110;
  40'd1582: rad_tmp = 24'b001011010010001101101110;
  40'd1583: rad_tmp = 24'b001011010010001101101110;
  40'd1584: rad_tmp = 24'b001011010011110100101011;
  40'd1585: rad_tmp = 24'b001011010011110100101011;
  40'd1586: rad_tmp = 24'b001011010011110100101011;
  40'd1587: rad_tmp = 24'b001011010011110100101011;
  40'd1588: rad_tmp = 24'b001011010011110100101011;
  40'd1589: rad_tmp = 24'b001011010011110100101011;
  40'd1590: rad_tmp = 24'b001011010011110100101011;
  40'd1591: rad_tmp = 24'b001011010011110100101011;
  40'd1592: rad_tmp = 24'b001011010011110100101011;
  40'd1593: rad_tmp = 24'b001011010011110100101011;
  40'd1594: rad_tmp = 24'b001011010011110100101011;
  40'd1595: rad_tmp = 24'b001011010011110100101011;
  40'd1596: rad_tmp = 24'b001011010011110100101011;
  40'd1597: rad_tmp = 24'b001011010011110100101011;
  40'd1598: rad_tmp = 24'b001011010011110100101011;
  40'd1599: rad_tmp = 24'b001011010011110100101011;
  40'd1600: rad_tmp = 24'b001011010011110100101011;
  40'd1601: rad_tmp = 24'b001011010011110100101011;
  40'd1602: rad_tmp = 24'b001011010011110100101011;
  40'd1603: rad_tmp = 24'b001011010011110100101011;
  40'd1604: rad_tmp = 24'b001011010011110100101011;
  40'd1605: rad_tmp = 24'b001011010011110100101011;
  40'd1606: rad_tmp = 24'b001011010011110100101011;
  40'd1607: rad_tmp = 24'b001011010011110100101011;
  40'd1608: rad_tmp = 24'b001011010011110100101011;
  40'd1609: rad_tmp = 24'b001011010011110100101011;
  40'd1610: rad_tmp = 24'b001011010011110100101011;
  40'd1611: rad_tmp = 24'b001011010011110100101011;
  40'd1612: rad_tmp = 24'b001011010011110100101011;
  40'd1613: rad_tmp = 24'b001011010011110100101011;
  40'd1614: rad_tmp = 24'b001011010011110100101011;
  40'd1615: rad_tmp = 24'b001011010011110100101011;
  40'd1616: rad_tmp = 24'b001011010101011011100111;
  40'd1617: rad_tmp = 24'b001011010101011011100111;
  40'd1618: rad_tmp = 24'b001011010101011011100111;
  40'd1619: rad_tmp = 24'b001011010101011011100111;
  40'd1620: rad_tmp = 24'b001011010101011011100111;
  40'd1621: rad_tmp = 24'b001011010101011011100111;
  40'd1622: rad_tmp = 24'b001011010101011011100111;
  40'd1623: rad_tmp = 24'b001011010101011011100111;
  40'd1624: rad_tmp = 24'b001011010101011011100111;
  40'd1625: rad_tmp = 24'b001011010101011011100111;
  40'd1626: rad_tmp = 24'b001011010101011011100111;
  40'd1627: rad_tmp = 24'b001011010101011011100111;
  40'd1628: rad_tmp = 24'b001011010101011011100111;
  40'd1629: rad_tmp = 24'b001011010101011011100111;
  40'd1630: rad_tmp = 24'b001011010101011011100111;
  40'd1631: rad_tmp = 24'b001011010101011011100111;
  40'd1632: rad_tmp = 24'b001011010101011011100111;
  40'd1633: rad_tmp = 24'b001011010101011011100111;
  40'd1634: rad_tmp = 24'b001011010101011011100111;
  40'd1635: rad_tmp = 24'b001011010101011011100111;
  40'd1636: rad_tmp = 24'b001011010101011011100111;
  40'd1637: rad_tmp = 24'b001011010101011011100111;
  40'd1638: rad_tmp = 24'b001011010101011011100111;
  40'd1639: rad_tmp = 24'b001011010101011011100111;
  40'd1640: rad_tmp = 24'b001011010101011011100111;
  40'd1641: rad_tmp = 24'b001011010101011011100111;
  40'd1642: rad_tmp = 24'b001011010101011011100111;
  40'd1643: rad_tmp = 24'b001011010101011011100111;
  40'd1644: rad_tmp = 24'b001011010101011011100111;
  40'd1645: rad_tmp = 24'b001011010101011011100111;
  40'd1646: rad_tmp = 24'b001011010101011011100111;
  40'd1647: rad_tmp = 24'b001011010101011011100111;
  40'd1648: rad_tmp = 24'b001011010101011011100111;
  40'd1649: rad_tmp = 24'b001011010101011011100111;
  40'd1650: rad_tmp = 24'b001011010111000010100100;
  40'd1651: rad_tmp = 24'b001011010111000010100100;
  40'd1652: rad_tmp = 24'b001011010111000010100100;
  40'd1653: rad_tmp = 24'b001011010111000010100100;
  40'd1654: rad_tmp = 24'b001011010111000010100100;
  40'd1655: rad_tmp = 24'b001011010111000010100100;
  40'd1656: rad_tmp = 24'b001011010111000010100100;
  40'd1657: rad_tmp = 24'b001011010111000010100100;
  40'd1658: rad_tmp = 24'b001011010111000010100100;
  40'd1659: rad_tmp = 24'b001011010111000010100100;
  40'd1660: rad_tmp = 24'b001011010111000010100100;
  40'd1661: rad_tmp = 24'b001011010111000010100100;
  40'd1662: rad_tmp = 24'b001011010111000010100100;
  40'd1663: rad_tmp = 24'b001011010111000010100100;
  40'd1664: rad_tmp = 24'b001011010111000010100100;
  40'd1665: rad_tmp = 24'b001011010111000010100100;
  40'd1666: rad_tmp = 24'b001011010111000010100100;
  40'd1667: rad_tmp = 24'b001011010111000010100100;
  40'd1668: rad_tmp = 24'b001011010111000010100100;
  40'd1669: rad_tmp = 24'b001011010111000010100100;
  40'd1670: rad_tmp = 24'b001011010111000010100100;
  40'd1671: rad_tmp = 24'b001011010111000010100100;
  40'd1672: rad_tmp = 24'b001011010111000010100100;
  40'd1673: rad_tmp = 24'b001011010111000010100100;
  40'd1674: rad_tmp = 24'b001011010111000010100100;
  40'd1675: rad_tmp = 24'b001011010111000010100100;
  40'd1676: rad_tmp = 24'b001011010111000010100100;
  40'd1677: rad_tmp = 24'b001011010111000010100100;
  40'd1678: rad_tmp = 24'b001011010111000010100100;
  40'd1679: rad_tmp = 24'b001011010111000010100100;
  40'd1680: rad_tmp = 24'b001011010111000010100100;
  40'd1681: rad_tmp = 24'b001011010111000010100100;
  40'd1682: rad_tmp = 24'b001011010111000010100100;
  40'd1683: rad_tmp = 24'b001011010111000010100100;
  40'd1684: rad_tmp = 24'b001011010111000010100100;
  40'd1685: rad_tmp = 24'b001011011000101001100000;
  40'd1686: rad_tmp = 24'b001011011000101001100000;
  40'd1687: rad_tmp = 24'b001011011000101001100000;
  40'd1688: rad_tmp = 24'b001011011000101001100000;
  40'd1689: rad_tmp = 24'b001011011000101001100000;
  40'd1690: rad_tmp = 24'b001011011000101001100000;
  40'd1691: rad_tmp = 24'b001011011000101001100000;
  40'd1692: rad_tmp = 24'b001011011000101001100000;
  40'd1693: rad_tmp = 24'b001011011000101001100000;
  40'd1694: rad_tmp = 24'b001011011000101001100000;
  40'd1695: rad_tmp = 24'b001011011000101001100000;
  40'd1696: rad_tmp = 24'b001011011000101001100000;
  40'd1697: rad_tmp = 24'b001011011000101001100000;
  40'd1698: rad_tmp = 24'b001011011000101001100000;
  40'd1699: rad_tmp = 24'b001011011000101001100000;
  40'd1700: rad_tmp = 24'b001011011000101001100000;
  40'd1701: rad_tmp = 24'b001011011000101001100000;
  40'd1702: rad_tmp = 24'b001011011000101001100000;
  40'd1703: rad_tmp = 24'b001011011000101001100000;
  40'd1704: rad_tmp = 24'b001011011000101001100000;
  40'd1705: rad_tmp = 24'b001011011000101001100000;
  40'd1706: rad_tmp = 24'b001011011000101001100000;
  40'd1707: rad_tmp = 24'b001011011000101001100000;
  40'd1708: rad_tmp = 24'b001011011000101001100000;
  40'd1709: rad_tmp = 24'b001011011000101001100000;
  40'd1710: rad_tmp = 24'b001011011000101001100000;
  40'd1711: rad_tmp = 24'b001011011000101001100000;
  40'd1712: rad_tmp = 24'b001011011000101001100000;
  40'd1713: rad_tmp = 24'b001011011000101001100000;
  40'd1714: rad_tmp = 24'b001011011000101001100000;
  40'd1715: rad_tmp = 24'b001011011000101001100000;
  40'd1716: rad_tmp = 24'b001011011000101001100000;
  40'd1717: rad_tmp = 24'b001011011000101001100000;
  40'd1718: rad_tmp = 24'b001011011000101001100000;
  40'd1719: rad_tmp = 24'b001011011000101001100000;
  40'd1720: rad_tmp = 24'b001011011000101001100000;
  40'd1721: rad_tmp = 24'b001011011010010000011100;
  40'd1722: rad_tmp = 24'b001011011010010000011100;
  40'd1723: rad_tmp = 24'b001011011010010000011100;
  40'd1724: rad_tmp = 24'b001011011010010000011100;
  40'd1725: rad_tmp = 24'b001011011010010000011100;
  40'd1726: rad_tmp = 24'b001011011010010000011100;
  40'd1727: rad_tmp = 24'b001011011010010000011100;
  40'd1728: rad_tmp = 24'b001011011010010000011100;
  40'd1729: rad_tmp = 24'b001011011010010000011100;
  40'd1730: rad_tmp = 24'b001011011010010000011100;
  40'd1731: rad_tmp = 24'b001011011010010000011100;
  40'd1732: rad_tmp = 24'b001011011010010000011100;
  40'd1733: rad_tmp = 24'b001011011010010000011100;
  40'd1734: rad_tmp = 24'b001011011010010000011100;
  40'd1735: rad_tmp = 24'b001011011010010000011100;
  40'd1736: rad_tmp = 24'b001011011010010000011100;
  40'd1737: rad_tmp = 24'b001011011010010000011100;
  40'd1738: rad_tmp = 24'b001011011010010000011100;
  40'd1739: rad_tmp = 24'b001011011010010000011100;
  40'd1740: rad_tmp = 24'b001011011010010000011100;
  40'd1741: rad_tmp = 24'b001011011010010000011100;
  40'd1742: rad_tmp = 24'b001011011010010000011100;
  40'd1743: rad_tmp = 24'b001011011010010000011100;
  40'd1744: rad_tmp = 24'b001011011010010000011100;
  40'd1745: rad_tmp = 24'b001011011010010000011100;
  40'd1746: rad_tmp = 24'b001011011010010000011100;
  40'd1747: rad_tmp = 24'b001011011010010000011100;
  40'd1748: rad_tmp = 24'b001011011010010000011100;
  40'd1749: rad_tmp = 24'b001011011010010000011100;
  40'd1750: rad_tmp = 24'b001011011010010000011100;
  40'd1751: rad_tmp = 24'b001011011010010000011100;
  40'd1752: rad_tmp = 24'b001011011010010000011100;
  40'd1753: rad_tmp = 24'b001011011010010000011100;
  40'd1754: rad_tmp = 24'b001011011010010000011100;
  40'd1755: rad_tmp = 24'b001011011010010000011100;
  40'd1756: rad_tmp = 24'b001011011010010000011100;
  40'd1757: rad_tmp = 24'b001011011010010000011100;
  40'd1758: rad_tmp = 24'b001011011010010000011100;
  40'd1759: rad_tmp = 24'b001011011011110111011001;
  40'd1760: rad_tmp = 24'b001011011011110111011001;
  40'd1761: rad_tmp = 24'b001011011011110111011001;
  40'd1762: rad_tmp = 24'b001011011011110111011001;
  40'd1763: rad_tmp = 24'b001011011011110111011001;
  40'd1764: rad_tmp = 24'b001011011011110111011001;
  40'd1765: rad_tmp = 24'b001011011011110111011001;
  40'd1766: rad_tmp = 24'b001011011011110111011001;
  40'd1767: rad_tmp = 24'b001011011011110111011001;
  40'd1768: rad_tmp = 24'b001011011011110111011001;
  40'd1769: rad_tmp = 24'b001011011011110111011001;
  40'd1770: rad_tmp = 24'b001011011011110111011001;
  40'd1771: rad_tmp = 24'b001011011011110111011001;
  40'd1772: rad_tmp = 24'b001011011011110111011001;
  40'd1773: rad_tmp = 24'b001011011011110111011001;
  40'd1774: rad_tmp = 24'b001011011011110111011001;
  40'd1775: rad_tmp = 24'b001011011011110111011001;
  40'd1776: rad_tmp = 24'b001011011011110111011001;
  40'd1777: rad_tmp = 24'b001011011011110111011001;
  40'd1778: rad_tmp = 24'b001011011011110111011001;
  40'd1779: rad_tmp = 24'b001011011011110111011001;
  40'd1780: rad_tmp = 24'b001011011011110111011001;
  40'd1781: rad_tmp = 24'b001011011011110111011001;
  40'd1782: rad_tmp = 24'b001011011011110111011001;
  40'd1783: rad_tmp = 24'b001011011011110111011001;
  40'd1784: rad_tmp = 24'b001011011011110111011001;
  40'd1785: rad_tmp = 24'b001011011011110111011001;
  40'd1786: rad_tmp = 24'b001011011011110111011001;
  40'd1787: rad_tmp = 24'b001011011011110111011001;
  40'd1788: rad_tmp = 24'b001011011011110111011001;
  40'd1789: rad_tmp = 24'b001011011011110111011001;
  40'd1790: rad_tmp = 24'b001011011011110111011001;
  40'd1791: rad_tmp = 24'b001011011011110111011001;
  40'd1792: rad_tmp = 24'b001011011011110111011001;
  40'd1793: rad_tmp = 24'b001011011011110111011001;
  40'd1794: rad_tmp = 24'b001011011011110111011001;
  40'd1795: rad_tmp = 24'b001011011011110111011001;
  40'd1796: rad_tmp = 24'b001011011011110111011001;
  40'd1797: rad_tmp = 24'b001011011011110111011001;
  40'd1798: rad_tmp = 24'b001011011011110111011001;
  40'd1799: rad_tmp = 24'b001011011101011110010101;
  40'd1800: rad_tmp = 24'b001011011101011110010101;
  40'd1801: rad_tmp = 24'b001011011101011110010101;
  40'd1802: rad_tmp = 24'b001011011101011110010101;
  40'd1803: rad_tmp = 24'b001011011101011110010101;
  40'd1804: rad_tmp = 24'b001011011101011110010101;
  40'd1805: rad_tmp = 24'b001011011101011110010101;
  40'd1806: rad_tmp = 24'b001011011101011110010101;
  40'd1807: rad_tmp = 24'b001011011101011110010101;
  40'd1808: rad_tmp = 24'b001011011101011110010101;
  40'd1809: rad_tmp = 24'b001011011101011110010101;
  40'd1810: rad_tmp = 24'b001011011101011110010101;
  40'd1811: rad_tmp = 24'b001011011101011110010101;
  40'd1812: rad_tmp = 24'b001011011101011110010101;
  40'd1813: rad_tmp = 24'b001011011101011110010101;
  40'd1814: rad_tmp = 24'b001011011101011110010101;
  40'd1815: rad_tmp = 24'b001011011101011110010101;
  40'd1816: rad_tmp = 24'b001011011101011110010101;
  40'd1817: rad_tmp = 24'b001011011101011110010101;
  40'd1818: rad_tmp = 24'b001011011101011110010101;
  40'd1819: rad_tmp = 24'b001011011101011110010101;
  40'd1820: rad_tmp = 24'b001011011101011110010101;
  40'd1821: rad_tmp = 24'b001011011101011110010101;
  40'd1822: rad_tmp = 24'b001011011101011110010101;
  40'd1823: rad_tmp = 24'b001011011101011110010101;
  40'd1824: rad_tmp = 24'b001011011101011110010101;
  40'd1825: rad_tmp = 24'b001011011101011110010101;
  40'd1826: rad_tmp = 24'b001011011101011110010101;
  40'd1827: rad_tmp = 24'b001011011101011110010101;
  40'd1828: rad_tmp = 24'b001011011101011110010101;
  40'd1829: rad_tmp = 24'b001011011101011110010101;
  40'd1830: rad_tmp = 24'b001011011101011110010101;
  40'd1831: rad_tmp = 24'b001011011101011110010101;
  40'd1832: rad_tmp = 24'b001011011101011110010101;
  40'd1833: rad_tmp = 24'b001011011101011110010101;
  40'd1834: rad_tmp = 24'b001011011101011110010101;
  40'd1835: rad_tmp = 24'b001011011101011110010101;
  40'd1836: rad_tmp = 24'b001011011101011110010101;
  40'd1837: rad_tmp = 24'b001011011101011110010101;
  40'd1838: rad_tmp = 24'b001011011101011110010101;
  40'd1839: rad_tmp = 24'b001011011101011110010101;
  40'd1840: rad_tmp = 24'b001011011111000101010010;
  40'd1841: rad_tmp = 24'b001011011111000101010010;
  40'd1842: rad_tmp = 24'b001011011111000101010010;
  40'd1843: rad_tmp = 24'b001011011111000101010010;
  40'd1844: rad_tmp = 24'b001011011111000101010010;
  40'd1845: rad_tmp = 24'b001011011111000101010010;
  40'd1846: rad_tmp = 24'b001011011111000101010010;
  40'd1847: rad_tmp = 24'b001011011111000101010010;
  40'd1848: rad_tmp = 24'b001011011111000101010010;
  40'd1849: rad_tmp = 24'b001011011111000101010010;
  40'd1850: rad_tmp = 24'b001011011111000101010010;
  40'd1851: rad_tmp = 24'b001011011111000101010010;
  40'd1852: rad_tmp = 24'b001011011111000101010010;
  40'd1853: rad_tmp = 24'b001011011111000101010010;
  40'd1854: rad_tmp = 24'b001011011111000101010010;
  40'd1855: rad_tmp = 24'b001011011111000101010010;
  40'd1856: rad_tmp = 24'b001011011111000101010010;
  40'd1857: rad_tmp = 24'b001011011111000101010010;
  40'd1858: rad_tmp = 24'b001011011111000101010010;
  40'd1859: rad_tmp = 24'b001011011111000101010010;
  40'd1860: rad_tmp = 24'b001011011111000101010010;
  40'd1861: rad_tmp = 24'b001011011111000101010010;
  40'd1862: rad_tmp = 24'b001011011111000101010010;
  40'd1863: rad_tmp = 24'b001011011111000101010010;
  40'd1864: rad_tmp = 24'b001011011111000101010010;
  40'd1865: rad_tmp = 24'b001011011111000101010010;
  40'd1866: rad_tmp = 24'b001011011111000101010010;
  40'd1867: rad_tmp = 24'b001011011111000101010010;
  40'd1868: rad_tmp = 24'b001011011111000101010010;
  40'd1869: rad_tmp = 24'b001011011111000101010010;
  40'd1870: rad_tmp = 24'b001011011111000101010010;
  40'd1871: rad_tmp = 24'b001011011111000101010010;
  40'd1872: rad_tmp = 24'b001011011111000101010010;
  40'd1873: rad_tmp = 24'b001011011111000101010010;
  40'd1874: rad_tmp = 24'b001011011111000101010010;
  40'd1875: rad_tmp = 24'b001011011111000101010010;
  40'd1876: rad_tmp = 24'b001011011111000101010010;
  40'd1877: rad_tmp = 24'b001011011111000101010010;
  40'd1878: rad_tmp = 24'b001011011111000101010010;
  40'd1879: rad_tmp = 24'b001011011111000101010010;
  40'd1880: rad_tmp = 24'b001011011111000101010010;
  40'd1881: rad_tmp = 24'b001011011111000101010010;
  40'd1882: rad_tmp = 24'b001011011111000101010010;
  40'd1883: rad_tmp = 24'b001011011111000101010010;
  40'd1884: rad_tmp = 24'b001011100000101100001110;
  40'd1885: rad_tmp = 24'b001011100000101100001110;
  40'd1886: rad_tmp = 24'b001011100000101100001110;
  40'd1887: rad_tmp = 24'b001011100000101100001110;
  40'd1888: rad_tmp = 24'b001011100000101100001110;
  40'd1889: rad_tmp = 24'b001011100000101100001110;
  40'd1890: rad_tmp = 24'b001011100000101100001110;
  40'd1891: rad_tmp = 24'b001011100000101100001110;
  40'd1892: rad_tmp = 24'b001011100000101100001110;
  40'd1893: rad_tmp = 24'b001011100000101100001110;
  40'd1894: rad_tmp = 24'b001011100000101100001110;
  40'd1895: rad_tmp = 24'b001011100000101100001110;
  40'd1896: rad_tmp = 24'b001011100000101100001110;
  40'd1897: rad_tmp = 24'b001011100000101100001110;
  40'd1898: rad_tmp = 24'b001011100000101100001110;
  40'd1899: rad_tmp = 24'b001011100000101100001110;
  40'd1900: rad_tmp = 24'b001011100000101100001110;
  40'd1901: rad_tmp = 24'b001011100000101100001110;
  40'd1902: rad_tmp = 24'b001011100000101100001110;
  40'd1903: rad_tmp = 24'b001011100000101100001110;
  40'd1904: rad_tmp = 24'b001011100000101100001110;
  40'd1905: rad_tmp = 24'b001011100000101100001110;
  40'd1906: rad_tmp = 24'b001011100000101100001110;
  40'd1907: rad_tmp = 24'b001011100000101100001110;
  40'd1908: rad_tmp = 24'b001011100000101100001110;
  40'd1909: rad_tmp = 24'b001011100000101100001110;
  40'd1910: rad_tmp = 24'b001011100000101100001110;
  40'd1911: rad_tmp = 24'b001011100000101100001110;
  40'd1912: rad_tmp = 24'b001011100000101100001110;
  40'd1913: rad_tmp = 24'b001011100000101100001110;
  40'd1914: rad_tmp = 24'b001011100000101100001110;
  40'd1915: rad_tmp = 24'b001011100000101100001110;
  40'd1916: rad_tmp = 24'b001011100000101100001110;
  40'd1917: rad_tmp = 24'b001011100000101100001110;
  40'd1918: rad_tmp = 24'b001011100000101100001110;
  40'd1919: rad_tmp = 24'b001011100000101100001110;
  40'd1920: rad_tmp = 24'b001011100000101100001110;
  40'd1921: rad_tmp = 24'b001011100000101100001110;
  40'd1922: rad_tmp = 24'b001011100000101100001110;
  40'd1923: rad_tmp = 24'b001011100000101100001110;
  40'd1924: rad_tmp = 24'b001011100000101100001110;
  40'd1925: rad_tmp = 24'b001011100000101100001110;
  40'd1926: rad_tmp = 24'b001011100000101100001110;
  40'd1927: rad_tmp = 24'b001011100000101100001110;
  40'd1928: rad_tmp = 24'b001011100000101100001110;
  40'd1929: rad_tmp = 24'b001011100010010011001010;
  40'd1930: rad_tmp = 24'b001011100010010011001010;
  40'd1931: rad_tmp = 24'b001011100010010011001010;
  40'd1932: rad_tmp = 24'b001011100010010011001010;
  40'd1933: rad_tmp = 24'b001011100010010011001010;
  40'd1934: rad_tmp = 24'b001011100010010011001010;
  40'd1935: rad_tmp = 24'b001011100010010011001010;
  40'd1936: rad_tmp = 24'b001011100010010011001010;
  40'd1937: rad_tmp = 24'b001011100010010011001010;
  40'd1938: rad_tmp = 24'b001011100010010011001010;
  40'd1939: rad_tmp = 24'b001011100010010011001010;
  40'd1940: rad_tmp = 24'b001011100010010011001010;
  40'd1941: rad_tmp = 24'b001011100010010011001010;
  40'd1942: rad_tmp = 24'b001011100010010011001010;
  40'd1943: rad_tmp = 24'b001011100010010011001010;
  40'd1944: rad_tmp = 24'b001011100010010011001010;
  40'd1945: rad_tmp = 24'b001011100010010011001010;
  40'd1946: rad_tmp = 24'b001011100010010011001010;
  40'd1947: rad_tmp = 24'b001011100010010011001010;
  40'd1948: rad_tmp = 24'b001011100010010011001010;
  40'd1949: rad_tmp = 24'b001011100010010011001010;
  40'd1950: rad_tmp = 24'b001011100010010011001010;
  40'd1951: rad_tmp = 24'b001011100010010011001010;
  40'd1952: rad_tmp = 24'b001011100010010011001010;
  40'd1953: rad_tmp = 24'b001011100010010011001010;
  40'd1954: rad_tmp = 24'b001011100010010011001010;
  40'd1955: rad_tmp = 24'b001011100010010011001010;
  40'd1956: rad_tmp = 24'b001011100010010011001010;
  40'd1957: rad_tmp = 24'b001011100010010011001010;
  40'd1958: rad_tmp = 24'b001011100010010011001010;
  40'd1959: rad_tmp = 24'b001011100010010011001010;
  40'd1960: rad_tmp = 24'b001011100010010011001010;
  40'd1961: rad_tmp = 24'b001011100010010011001010;
  40'd1962: rad_tmp = 24'b001011100010010011001010;
  40'd1963: rad_tmp = 24'b001011100010010011001010;
  40'd1964: rad_tmp = 24'b001011100010010011001010;
  40'd1965: rad_tmp = 24'b001011100010010011001010;
  40'd1966: rad_tmp = 24'b001011100010010011001010;
  40'd1967: rad_tmp = 24'b001011100010010011001010;
  40'd1968: rad_tmp = 24'b001011100010010011001010;
  40'd1969: rad_tmp = 24'b001011100010010011001010;
  40'd1970: rad_tmp = 24'b001011100010010011001010;
  40'd1971: rad_tmp = 24'b001011100010010011001010;
  40'd1972: rad_tmp = 24'b001011100010010011001010;
  40'd1973: rad_tmp = 24'b001011100010010011001010;
  40'd1974: rad_tmp = 24'b001011100010010011001010;
  40'd1975: rad_tmp = 24'b001011100010010011001010;
  40'd1976: rad_tmp = 24'b001011100011111010000111;
  40'd1977: rad_tmp = 24'b001011100011111010000111;
  40'd1978: rad_tmp = 24'b001011100011111010000111;
  40'd1979: rad_tmp = 24'b001011100011111010000111;
  40'd1980: rad_tmp = 24'b001011100011111010000111;
  40'd1981: rad_tmp = 24'b001011100011111010000111;
  40'd1982: rad_tmp = 24'b001011100011111010000111;
  40'd1983: rad_tmp = 24'b001011100011111010000111;
  40'd1984: rad_tmp = 24'b001011100011111010000111;
  40'd1985: rad_tmp = 24'b001011100011111010000111;
  40'd1986: rad_tmp = 24'b001011100011111010000111;
  40'd1987: rad_tmp = 24'b001011100011111010000111;
  40'd1988: rad_tmp = 24'b001011100011111010000111;
  40'd1989: rad_tmp = 24'b001011100011111010000111;
  40'd1990: rad_tmp = 24'b001011100011111010000111;
  40'd1991: rad_tmp = 24'b001011100011111010000111;
  40'd1992: rad_tmp = 24'b001011100011111010000111;
  40'd1993: rad_tmp = 24'b001011100011111010000111;
  40'd1994: rad_tmp = 24'b001011100011111010000111;
  40'd1995: rad_tmp = 24'b001011100011111010000111;
  40'd1996: rad_tmp = 24'b001011100011111010000111;
  40'd1997: rad_tmp = 24'b001011100011111010000111;
  40'd1998: rad_tmp = 24'b001011100011111010000111;
  40'd1999: rad_tmp = 24'b001011100011111010000111;
  40'd2000: rad_tmp = 24'b001011100011111010000111;
  40'd2001: rad_tmp = 23'b001011100011111010000111;
  40'd2002: rad_tmp = 23'b001011100011111010000111;
  40'd2003: rad_tmp = 23'b001011100011111010000111;
  40'd2004: rad_tmp = 23'b001011100011111010000111;
  40'd2005: rad_tmp = 23'b001011100011111010000111;
  40'd2006: rad_tmp = 23'b001011100011111010000111;
  40'd2007: rad_tmp = 23'b001011100011111010000111;
  40'd2008: rad_tmp = 23'b001011100011111010000111;
  40'd2009: rad_tmp = 23'b001011100011111010000111;
  40'd2010: rad_tmp = 23'b001011100011111010000111;
  40'd2011: rad_tmp = 23'b001011100011111010000111;
  40'd2012: rad_tmp = 23'b001011100011111010000111;
  40'd2013: rad_tmp = 23'b001011100011111010000111;
  40'd2014: rad_tmp = 23'b001011100011111010000111;
  40'd2015: rad_tmp = 23'b001011100011111010000111;
  40'd2016: rad_tmp = 23'b001011100011111010000111;
  40'd2017: rad_tmp = 23'b001011100011111010000111;
  40'd2018: rad_tmp = 23'b001011100011111010000111;
  40'd2019: rad_tmp = 23'b001011100011111010000111;
  40'd2020: rad_tmp = 23'b001011100011111010000111;
  40'd2021: rad_tmp = 23'b001011100011111010000111;
  40'd2022: rad_tmp = 23'b001011100011111010000111;
  40'd2023: rad_tmp = 23'b001011100011111010000111;
  40'd2024: rad_tmp = 23'b001011100011111010000111;
  40'd2025: rad_tmp = 23'b001011100011111010000111;
  40'd2026: rad_tmp = 23'b001011100101100001000011;
  40'd2027: rad_tmp = 23'b001011100101100001000011;
  40'd2028: rad_tmp = 23'b001011100101100001000011;
  40'd2029: rad_tmp = 23'b001011100101100001000011;
  40'd2030: rad_tmp = 23'b001011100101100001000011;
  40'd2031: rad_tmp = 23'b001011100101100001000011;
  40'd2032: rad_tmp = 23'b001011100101100001000011;
  40'd2033: rad_tmp = 23'b001011100101100001000011;
  40'd2034: rad_tmp = 23'b001011100101100001000011;
  40'd2035: rad_tmp = 23'b001011100101100001000011;
  40'd2036: rad_tmp = 23'b001011100101100001000011;
  40'd2037: rad_tmp = 23'b001011100101100001000011;
  40'd2038: rad_tmp = 23'b001011100101100001000011;
  40'd2039: rad_tmp = 23'b001011100101100001000011;
  40'd2040: rad_tmp = 23'b001011100101100001000011;
  40'd2041: rad_tmp = 23'b001011100101100001000011;
  40'd2042: rad_tmp = 23'b001011100101100001000011;
  40'd2043: rad_tmp = 23'b001011100101100001000011;
  40'd2044: rad_tmp = 23'b001011100101100001000011;
  40'd2045: rad_tmp = 23'b001011100101100001000011;
  40'd2046: rad_tmp = 23'b001011100101100001000011;
  40'd2047: rad_tmp = 23'b001011100101100001000011;
endcase
end
end
endmodule
