`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2018/08/18 12:06:47
// Design Name:
// Module Name: CAL_Module
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module CAL_Module(
  input wire clk,
  input wire rst,
  input wire input_valid,
  input wire [576 : 1] wm_data,
  input wire [576 : 1] i_data,
  output wire [576 : 1] o_data
    );
    
    
    wire  [18:1] i_imag_Y1 [8:1];
    wire  [18:1] i_imag_Y2 [8:1];
    wire  [18:1] i_imag_Y3 [8:1];
    wire  [18:1] i_imag_U1 [8:1];
    wire  [18:1] i_imag_U2 [8:1];
    wire  [18:1] i_imag_U3 [8:1];
    wire  [18:1] i_imag_V1 [8:1];
    wire  [18:1] i_imag_V2 [8:1];
    wire  [18:1] i_imag_V3 [8:1];
    wire  [576:1]data          ;
    wire  signed [19:1] o_imag_Y1 [8:1];
    wire  signed [19:1] o_imag_Y2 [8:1];
    wire  signed [19:1] o_imag_Y3 [8:1];
    wire  signed [19:1] o_imag_U1 [8:1];
    wire  signed [19:1] o_imag_U2 [8:1];
    wire  signed [19:1] o_imag_U3 [8:1];
    wire  signed [19:1] o_imag_V1 [8:1];
    wire  signed [19:1] o_imag_V2 [8:1];
    wire  signed [19:1] o_imag_V3 [8:1];
    
    wire  [29:1] o_imag_R1 [8:1];
    wire  [29:1] o_imag_R2 [8:1];
    wire  [29:1] o_imag_R3 [8:1];
    wire  [29:1] o_imag_G1 [8:1];
    wire  [29:1] o_imag_G2 [8:1];
    wire  [29:1] o_imag_G3 [8:1];
    wire  [29:1] o_imag_B1 [8:1];
    wire  [29:1] o_imag_B2 [8:1];
    wire  [29:1] o_imag_B3 [8:1];
    
    wire  [8:1] o_imag_R1_f [8:1];
    wire  [8:1] o_imag_R2_f [8:1];
    wire  [8:1] o_imag_R3_f [8:1];
    wire  [8:1] o_imag_G1_f [8:1];
    wire  [8:1] o_imag_G2_f [8:1];
    wire  [8:1] o_imag_G3_f [8:1];
    wire  [8:1] o_imag_B1_f [8:1];
    wire  [8:1] o_imag_B2_f [8:1];
    wire  [8:1] o_imag_B3_f [8:1];
    
     assign o_imag_R1_f[1] = o_imag_R1[1][28:21] + o_imag_R1[1][20];
     assign o_imag_R1_f[2] = o_imag_R1[2][28:21] + o_imag_R1[2][20];
     assign o_imag_R1_f[3] = o_imag_R1[3][28:21] + o_imag_R1[3][20];
     assign o_imag_R1_f[4] = o_imag_R1[4][28:21] + o_imag_R1[4][20];
     assign o_imag_R1_f[5] = o_imag_R1[5][28:21] + o_imag_R1[5][20];
     assign o_imag_R1_f[6] = o_imag_R1[6][28:21] + o_imag_R1[6][20];
     assign o_imag_R1_f[7] = o_imag_R1[7][28:21] + o_imag_R1[7][20];
     assign o_imag_R1_f[8] = o_imag_R1[8][28:21] + o_imag_R1[8][20];
     //R2          R=_f o_ =        R= o_[28:21] +        R= o_[20];
     assign o_imag_R2_f[1] = o_imag_R2[1][28:21] + o_imag_R2[1][20];
     assign o_imag_R2_f[2] = o_imag_R2[2][28:21] + o_imag_R2[2][20];
     assign o_imag_R2_f[3] = o_imag_R2[3][28:21] + o_imag_R2[3][20];
     assign o_imag_R2_f[4] = o_imag_R2[4][28:21] + o_imag_R2[4][20];
     assign o_imag_R2_f[5] = o_imag_R2[5][28:21] + o_imag_R2[5][20];
     assign o_imag_R2_f[6] = o_imag_R2[6][28:21] + o_imag_R2[6][20];
     assign o_imag_R2_f[7] = o_imag_R2[7][28:21] + o_imag_R2[7][20];
     assign o_imag_R2_f[8] = o_imag_R2[8][28:21] + o_imag_R2[8][20];
      //R3         R _f= o =        R = o[28:21] +        R = o[20];
     assign o_imag_R3_f[1] = o_imag_R3[1][28:21] + o_imag_R3[1][20];
     assign o_imag_R3_f[2] = o_imag_R3[2][28:21] + o_imag_R3[2][20];
     assign o_imag_R3_f[3] = o_imag_R3[3][28:21] + o_imag_R3[3][20];
     assign o_imag_R3_f[4] = o_imag_R3[4][28:21] + o_imag_R3[4][20];
     assign o_imag_R3_f[5] = o_imag_R3[5][28:21] + o_imag_R3[5][20];
     assign o_imag_R3_f[6] = o_imag_R3[6][28:21] + o_imag_R3[6][20];
     assign o_imag_R3_f[7] = o_imag_R3[7][28:21] + o_imag_R3[7][20];
     assign o_imag_R3_f[8] = o_imag_R3[8][28:21] + o_imag_R3[8][20];
     //   G=Y-0.34414_f*(U = Y-0.34414*(U[28:21] + Y-0.34414*(U[20];
     //G1            _f    =             [28:21] +             [20];
     assign o_imag_G1_f[1] = o_imag_G1[1][28:21] + o_imag_G1[1][20];
     assign o_imag_G1_f[2] = o_imag_G1[2][28:21] + o_imag_G1[2][20];
     assign o_imag_G1_f[3] = o_imag_G1[3][28:21] + o_imag_G1[3][20];
     assign o_imag_G1_f[4] = o_imag_G1[4][28:21] + o_imag_G1[4][20];
     assign o_imag_G1_f[5] = o_imag_G1[5][28:21] + o_imag_G1[5][20];
     assign o_imag_G1_f[6] = o_imag_G1[6][28:21] + o_imag_G1[6][20];
     assign o_imag_G1_f[7] = o_imag_G1[7][28:21] + o_imag_G1[7][20];
     assign o_imag_G1_f[8] = o_imag_G1[8][28:21] + o_imag_G1[8][20];
      //G2   G     G _f= o =  G     G = o[28:21] +  G     G = o[20];
     assign o_imag_G2_f[1] = o_imag_G2[1][28:21] + o_imag_G2[1][20];
     assign o_imag_G2_f[2] = o_imag_G2[2][28:21] + o_imag_G2[2][20];
     assign o_imag_G2_f[3] = o_imag_G2[3][28:21] + o_imag_G2[3][20];
     assign o_imag_G2_f[4] = o_imag_G2[4][28:21] + o_imag_G2[4][20];
     assign o_imag_G2_f[5] = o_imag_G2[5][28:21] + o_imag_G2[5][20];
     assign o_imag_G2_f[6] = o_imag_G2[6][28:21] + o_imag_G2[6][20];
     assign o_imag_G2_f[7] = o_imag_G2[7][28:21] + o_imag_G2[7][20];
     assign o_imag_G2_f[8] = o_imag_G2[8][28:21] + o_imag_G2[8][20];
     //G3   G      G=_f o_ = G      G= o_[28:21] + G      G= o_[20];
     assign o_imag_G3_f[1] = o_imag_G3[1][28:21] + o_imag_G3[1][20];
     assign o_imag_G3_f[2] = o_imag_G3[2][28:21] + o_imag_G3[2][20];
     assign o_imag_G3_f[3] = o_imag_G3[3][28:21] + o_imag_G3[3][20];
     assign o_imag_G3_f[4] = o_imag_G3[4][28:21] + o_imag_G3[4][20];
     assign o_imag_G3_f[5] = o_imag_G3[5][28:21] + o_imag_G3[5][20];
     assign o_imag_G3_f[6] = o_imag_G3[6][28:21] + o_imag_G3[6][20];
     assign o_imag_G3_f[7] = o_imag_G3[7][28:21] + o_imag_G3[7][20];
     assign o_imag_G3_f[8] = o_imag_G3[8][28:21] + o_imag_G3[8][20];
     //   B=Y+1.772G(_fU-1   Y+1.772G(U-1[28:21] + Y+1.772G(U-1[20];
     //R1            _f                  [28:21] +             [20];
     assign o_imag_B1_f[1] = o_imag_B1[1][28:21] + o_imag_B1[1][20];
     assign o_imag_B1_f[2] = o_imag_B1[2][28:21] + o_imag_B1[2][20];
     assign o_imag_B1_f[3] = o_imag_B1[3][28:21] + o_imag_B1[3][20];
     assign o_imag_B1_f[4] = o_imag_B1[4][28:21] + o_imag_B1[4][20];
     assign o_imag_B1_f[5] = o_imag_B1[5][28:21] + o_imag_B1[5][20];
     assign o_imag_B1_f[6] = o_imag_B1[6][28:21] + o_imag_B1[6][20];
     assign o_imag_B1_f[7] = o_imag_B1[7][28:21] + o_imag_B1[7][20];
     assign o_imag_B1_f[8] = o_imag_B1[8][28:21] + o_imag_B1[8][20];
     //R2   B      B=_f o_ = B      B= o_[28:21] + B      B= o_[20];
     assign o_imag_B2_f[1] = o_imag_B2[1][28:21] + o_imag_B2[1][20];
     assign o_imag_B2_f[2] = o_imag_B2[2][28:21] + o_imag_B2[2][20];
     assign o_imag_B2_f[3] = o_imag_B2[3][28:21] + o_imag_B2[3][20];
     assign o_imag_B2_f[4] = o_imag_B2[4][28:21] + o_imag_B2[4][20];
     assign o_imag_B2_f[5] = o_imag_B2[5][28:21] + o_imag_B2[5][20];
     assign o_imag_B2_f[6] = o_imag_B2[6][28:21] + o_imag_B2[6][20];
     assign o_imag_B2_f[7] = o_imag_B2[7][28:21] + o_imag_B2[7][20];
     assign o_imag_B2_f[8] = o_imag_B2[8][28:21] + o_imag_B2[8][20];
      //R3   B     B _f= o =  B     B = o[28:21] +  B     B = o[20];
     assign o_imag_B3_f[1] = o_imag_B3[1][28:21] + o_imag_B3[1][20];
     assign o_imag_B3_f[2] = o_imag_B3[2][28:21] + o_imag_B3[2][20];
     assign o_imag_B3_f[3] = o_imag_B3[3][28:21] + o_imag_B3[3][20];
     assign o_imag_B3_f[4] = o_imag_B3[4][28:21] + o_imag_B3[4][20];
     assign o_imag_B3_f[5] = o_imag_B3[5][28:21] + o_imag_B3[5][20];
     assign o_imag_B3_f[6] = o_imag_B3[6][28:21] + o_imag_B3[6][20];
     assign o_imag_B3_f[7] = o_imag_B3[7][28:21] + o_imag_B3[7][20];
     assign o_imag_B3_f[8] = o_imag_B3[8][28:21] + o_imag_B3[8][20];
     
     
    assign o_imag_Y1[1][19] = 1'b0;
    assign o_imag_Y1[2][19] = 1'b0;
    assign o_imag_Y1[3][19] = 1'b0;
    assign o_imag_Y1[4][19] = 1'b0;
    assign o_imag_Y1[5][19] = 1'b0;
    assign o_imag_Y1[6][19] = 1'b0;
    assign o_imag_Y1[7][19] = 1'b0;
    assign o_imag_Y1[8][19] = 1'b0;
    //R2          Y= o_[19]im 1'b0;
    assign o_imag_Y2[1][19] = 1'b0;
    assign o_imag_Y2[2][19] = 1'b0;
    assign o_imag_Y2[3][19] = 1'b0;
    assign o_imag_Y2[4][19] = 1'b0;
    assign o_imag_Y2[5][19] = 1'b0;
    assign o_imag_Y2[6][19] = 1'b0;
    assign o_imag_Y2[7][19] = 1'b0;
    assign o_imag_Y2[8][19] = 1'b0;
     //R3         Y = o[19]_i 1'b0;
    assign o_imag_Y3[1][19] = 1'b0;
    assign o_imag_Y3[2][19] = 1'b0;
    assign o_imag_Y3[3][19] = 1'b0;
    assign o_imag_Y3[4][19] = 1'b0;
    assign o_imag_Y3[5][19] = 1'b0;
    assign o_imag_Y3[6][19] = 1'b0;
    assign o_imag_Y3[7][19] = 1'b0;
    assign o_imag_Y3[8][19] = 1'b0;
    //   G=Y-0.34414*(U[19]-1 1'b0;
    //G1               [19]   1'b0;
    assign o_imag_U1[1][19] = 1'b0;
    assign o_imag_U1[2][19] = 1'b0;
    assign o_imag_U1[3][19] = 1'b0;
    assign o_imag_U1[4][19] = 1'b0;
    assign o_imag_U1[5][19] = 1'b0;
    assign o_imag_U1[6][19] = 1'b0;
    assign o_imag_U1[7][19] = 1'b0;
    assign o_imag_U1[8][19] = 1'b0;
     //G2   G     U = o[19]_i 1'b0;
    assign o_imag_U2[1][19] = 1'b0;
    assign o_imag_U2[2][19] = 1'b0;
    assign o_imag_U2[3][19] = 1'b0;
    assign o_imag_U2[4][19] = 1'b0;
    assign o_imag_U2[5][19] = 1'b0;
    assign o_imag_U2[6][19] = 1'b0;
    assign o_imag_U2[7][19] = 1'b0;
    assign o_imag_U2[8][19] = 1'b0;
    //G3   G      U= o_[19]im 1'b0;
    assign o_imag_U3[1][19] = 1'b0;
    assign o_imag_U3[2][19] = 1'b0;
    assign o_imag_U3[3][19] = 1'b0;
    assign o_imag_U3[4][19] = 1'b0;
    assign o_imag_U3[5][19] = 1'b0;
    assign o_imag_U3[6][19] = 1'b0;
    assign o_imag_U3[7][19] = 1'b0;
    assign o_imag_U3[8][19] = 1'b0;
    //   B=Y+1.772*(U-1[19]28 1'b0;
    //R1               [19]   1'b0;
    assign o_imag_V1[1][19] = 1'b0;
    assign o_imag_V1[2][19] = 1'b0;
    assign o_imag_V1[3][19] = 1'b0;
    assign o_imag_V1[4][19] = 1'b0;
    assign o_imag_V1[5][19] = 1'b0;
    assign o_imag_V1[6][19] = 1'b0;
    assign o_imag_V1[7][19] = 1'b0;
    assign o_imag_V1[8][19] = 1'b0;
    //R2   B      V= o_[19]im 1'b0;
    assign o_imag_V2[1][19] = 1'b0;
    assign o_imag_V2[2][19] = 1'b0;
    assign o_imag_V2[3][19] = 1'b0;
    assign o_imag_V2[4][19] = 1'b0;
    assign o_imag_V2[5][19] = 1'b0;
    assign o_imag_V2[6][19] = 1'b0;
    assign o_imag_V2[7][19] = 1'b0;
    assign o_imag_V2[8][19] = 1'b0;
     //R3   B     V = o[19]_i 1'b0;
    assign o_imag_V3[1][19] = 1'b0;
    assign o_imag_V3[2][19] = 1'b0;
    assign o_imag_V3[3][19] = 1'b0;
    assign o_imag_V3[4][19] = 1'b0;
    assign o_imag_V3[5][19] = 1'b0;
    assign o_imag_V3[6][19] = 1'b0;
    assign o_imag_V3[7][19] = 1'b0;
    assign o_imag_V3[8][19] = 1'b0;
  




    reg [30:1] cnt ;
    reg [30:1] cnt_cycle;
    reg [10:0] cnt_cycle_l;
    reg [18:1] wm;
    reg [18:1] watermark [2222:0];
    
    
    always@(posedge clk) begin
      if(rst == 1) begin
        cnt         <= 0;
        cnt_cycle   <= 0;
        cnt_cycle_l <= 0;
        
        watermark[0] <= 18'b111111111111111111;
        watermark[1] <= 18'b111111111111111111;
        watermark[2] <= 18'b111111111111111111;
        watermark[3] <= 18'b111111111111111111;
        watermark[4] <= 18'b111111111111111111;
        watermark[5] <= 18'b111111111111111111;
        watermark[6] <= 18'b111111111111111111;
        watermark[7] <= 18'b111111111111111111;
        watermark[8] <= 18'b111111111111111111;
        watermark[9] <= 18'b111111111111111111;
        watermark[10] <= 18'b111111111111111111;
        watermark[11] <= 18'b111111111111111111;
        watermark[12] <= 18'b111111111111111111;
        watermark[13] <= 18'b111111111111111111;
        watermark[14] <= 18'b111111111111111111;
        watermark[15] <= 18'b111111111111111111;
        watermark[16] <= 18'b111111111111111111;
        watermark[17] <= 18'b111111111111111111;
        watermark[18] <= 18'b111111111111111111;
        watermark[19] <= 18'b111111111111111111;
        watermark[20] <= 18'b111111111111111111;
        watermark[21] <= 18'b111111111111111111;
        watermark[22] <= 18'b111111111111111111;
        watermark[23] <= 18'b111111111111111111;
        watermark[24] <= 18'b111111111111111111;
        watermark[25] <= 18'b111111111111111111;
        watermark[26] <= 18'b111111111111111111;
        watermark[27] <= 18'b111111111111111111;
        watermark[28] <= 18'b111111111111111111;
        watermark[29] <= 18'b111111111111111111;
        watermark[30] <= 18'b111111111111111111;
        watermark[31] <= 18'b111111111111111111;
        watermark[32] <= 18'b111111111111111111;
        watermark[33] <= 18'b111111111111111111;
        watermark[34] <= 18'b111111111111111111;
        watermark[35] <= 18'b111111111111111111;
        watermark[36] <= 18'b111111111111111111;
        watermark[37] <= 18'b111111111111111111;
        watermark[38] <= 18'b111111111111111111;
        watermark[39] <= 18'b111111111111111111;
        watermark[40] <= 18'b111111111111111111;
        watermark[41] <= 18'b111111111111111111;
        watermark[42] <= 18'b111111111111111111;
        watermark[43] <= 18'b111111111111111111;
        watermark[44] <= 18'b111111111111111111;
        watermark[45] <= 18'b111111111111111111;
        watermark[46] <= 18'b111111111111111111;
        watermark[47] <= 18'b111111111111111111;
        watermark[48] <= 18'b111111111111111111;
        watermark[49] <= 18'b111111111111111111;
        watermark[50] <= 18'b111111111111111111;
        watermark[51] <= 18'b111111111111111111;
        watermark[52] <= 18'b111111111111111111;
        watermark[53] <= 18'b111111111111111111;
        watermark[54] <= 18'b111111111111111111;
        watermark[55] <= 18'b111111111111111111;
        watermark[56] <= 18'b111111111111111111;
        watermark[57] <= 18'b111111111111111111;
        watermark[58] <= 18'b111111111111111111;
        watermark[59] <= 18'b111111111111111111;
        watermark[60] <= 18'b111111111111111111;
        watermark[61] <= 18'b111111111111111111;
        watermark[62] <= 18'b111111111111111111;
        watermark[63] <= 18'b111111111111111111;
        watermark[64] <= 18'b111111111111111111;
        watermark[65] <= 18'b111111111111111111;
        watermark[66] <= 18'b111111111111111111;
        watermark[67] <= 18'b111111111111111111;
        watermark[68] <= 18'b111111111111111111;
        watermark[69] <= 18'b111111111111111111;
        watermark[70] <= 18'b111111111111111111;
        watermark[71] <= 18'b111111111111111111;
        watermark[72] <= 18'b111111111111111111;
        watermark[73] <= 18'b111111111111111111;
        watermark[74] <= 18'b111111111111111111;
        watermark[75] <= 18'b111111111111111111;
        watermark[76] <= 18'b111111111111111111;
        watermark[77] <= 18'b111111111111111111;
        watermark[78] <= 18'b111111111111111111;
        watermark[79] <= 18'b111111111111111111;
        watermark[80] <= 18'b111111111111111111;
        watermark[81] <= 18'b111111111111111111;
        watermark[82] <= 18'b111111111111111111;
        watermark[83] <= 18'b111111111111111111;
        watermark[84] <= 18'b111111111111111111;
        watermark[85] <= 18'b111111111111111111;
        watermark[86] <= 18'b111111111111111111;
        watermark[87] <= 18'b111111111111111111;
        watermark[88] <= 18'b111111111111111111;
        watermark[89] <= 18'b111111111111111111;
        watermark[90] <= 18'b111111111111111111;
        watermark[91] <= 18'b111111111111111111;
        watermark[92] <= 18'b111111111111111111;
        watermark[93] <= 18'b111111111111111111;
        watermark[94] <= 18'b111111111111111111;
        watermark[95] <= 18'b111111111111111111;
        watermark[96] <= 18'b111111111111111111;
        watermark[97] <= 18'b111111111111111111;
        watermark[98] <= 18'b111111111111111111;
        watermark[99] <= 18'b111111111111111111;
        watermark[100] <= 18'b111111111111111111;
        watermark[101] <= 18'b111111111111111111;
        watermark[102] <= 18'b111111111111111111;
        watermark[103] <= 18'b111111111111111111;
        watermark[104] <= 18'b111111111111111111;
        watermark[105] <= 18'b111111111111111111;
        watermark[106] <= 18'b111111111111111111;
        watermark[107] <= 18'b111111111111111111;
        watermark[108] <= 18'b111111111111111111;
        watermark[109] <= 18'b111111111111111111;
        watermark[110] <= 18'b111111111111111111;
        watermark[111] <= 18'b111111111111111111;
        watermark[112] <= 18'b111111111111111111;
        watermark[113] <= 18'b111111111111111111;
        watermark[114] <= 18'b111111111111111111;
        watermark[115] <= 18'b111111111111111111;
        watermark[116] <= 18'b111111111111111111;
        watermark[117] <= 18'b111111111111111111;
        watermark[118] <= 18'b111111111111111111;
        watermark[119] <= 18'b111111111111111111;
        watermark[120] <= 18'b111111111111111111;
        watermark[121] <= 18'b111111111111111111;
        watermark[122] <= 18'b111111111111111111;
        watermark[123] <= 18'b111111111111111111;
        watermark[124] <= 18'b111111111111111111;
        watermark[125] <= 18'b111111111111111111;
        watermark[126] <= 18'b111111111111111111;
        watermark[127] <= 18'b111111111111111111;
        watermark[128] <= 18'b111111111111111111;
        watermark[129] <= 18'b111111111111111111;
        watermark[130] <= 18'b111111111111111111;
        watermark[131] <= 18'b111111111111111111;
        watermark[132] <= 18'b111111111111111111;
        watermark[133] <= 18'b111111111111111111;
        watermark[134] <= 18'b111111111111111111;
        watermark[135] <= 18'b111111111111111111;
        watermark[136] <= 18'b111111111111111111;
        watermark[137] <= 18'b111111111111111111;
        watermark[138] <= 18'b111111111111111111;
        watermark[139] <= 18'b111111111111111111;
        watermark[140] <= 18'b111111111111111111;
        watermark[141] <= 18'b111111111111111111;
        watermark[142] <= 18'b111111111111111111;
        watermark[143] <= 18'b111111111111111111;
        watermark[144] <= 18'b111111111111111111;
        watermark[145] <= 18'b111111111111111111;
        watermark[146] <= 18'b111111111111111111;
        watermark[147] <= 18'b111111111111111111;
        watermark[148] <= 18'b111111111111111111;
        watermark[149] <= 18'b111111111111111111;
        watermark[150] <= 18'b111111111111111111;
        watermark[151] <= 18'b111111111111111111;
        watermark[152] <= 18'b111111111111111111;
        watermark[153] <= 18'b111111111111111111;
        watermark[154] <= 18'b111111111111111111;
        watermark[155] <= 18'b111111111111111111;
        watermark[156] <= 18'b111111111111111111;
        watermark[157] <= 18'b111111111111111111;
        watermark[158] <= 18'b111111111111111111;
        watermark[159] <= 18'b111111111111111111;
        watermark[160] <= 18'b111111111111111111;
        watermark[161] <= 18'b111111111111111111;
        watermark[162] <= 18'b111111111111111111;
        watermark[163] <= 18'b111111111111111111;
        watermark[164] <= 18'b111111111111111111;
        watermark[165] <= 18'b111111111111111111;
        watermark[166] <= 18'b111111111111111111;
        watermark[167] <= 18'b111111111111111111;
        watermark[168] <= 18'b111111111111111111;
        watermark[169] <= 18'b111111111111111111;
        watermark[170] <= 18'b111111111111111111;
        watermark[171] <= 18'b111111111111111111;
        watermark[172] <= 18'b111111111111111111;
        watermark[173] <= 18'b111111111111111111;
        watermark[174] <= 18'b111111111111111111;
        watermark[175] <= 18'b111111111111111111;
        watermark[176] <= 18'b111111111111111111;
        watermark[177] <= 18'b111111111111111111;
        watermark[178] <= 18'b111111111111111111;
        watermark[179] <= 18'b111111111111111111;
        watermark[180] <= 18'b111111111111111111;
        watermark[181] <= 18'b111111111111111111;
        watermark[182] <= 18'b111111111111111111;
        watermark[183] <= 18'b111111111111111111;
        watermark[184] <= 18'b111111111111111111;
        watermark[185] <= 18'b111111111111111111;
        watermark[186] <= 18'b111111111111111111;
        watermark[187] <= 18'b111111111111111111;
        watermark[188] <= 18'b111111111111111111;
        watermark[189] <= 18'b111111111111111111;
        watermark[190] <= 18'b111111111111111111;
        watermark[191] <= 18'b111111111111111111;
        watermark[192] <= 18'b111111111111111111;
        watermark[193] <= 18'b111111111111111111;
        watermark[194] <= 18'b111111111111111111;
        watermark[195] <= 18'b111111111111111111;
        watermark[196] <= 18'b111111111111111111;
        watermark[197] <= 18'b111111111111111111;
        watermark[198] <= 18'b111111111111111111;
        watermark[199] <= 18'b111111111111111111;
        watermark[200] <= 18'b111111111111111111;
        watermark[201] <= 18'b111111111111111111;
        watermark[202] <= 18'b111111111111111111;
        watermark[203] <= 18'b111111111111111111;
        watermark[204] <= 18'b111111111111111111;
        watermark[205] <= 18'b111111111111111111;
        watermark[206] <= 18'b111111111111111111;
        watermark[207] <= 18'b111111111111111111;
        watermark[208] <= 18'b111111111111111111;
        watermark[209] <= 18'b111111111111111111;
        watermark[210] <= 18'b111111111111111111;
        watermark[211] <= 18'b111111111111111111;
        watermark[212] <= 18'b111111111111111111;
        watermark[213] <= 18'b111111111111111111;
        watermark[214] <= 18'b111111111111111111;
        watermark[215] <= 18'b111111111111111111;
        watermark[216] <= 18'b111111111111111111;
        watermark[217] <= 18'b111111111111111111;
        watermark[218] <= 18'b111111111111111111;
        watermark[219] <= 18'b111111111111111111;
        watermark[220] <= 18'b111111111111111111;
        watermark[221] <= 18'b111111111111111111;
        watermark[222] <= 18'b111111111111111111;
        watermark[223] <= 18'b111111111111111111;
        watermark[224] <= 18'b111111111111111111;
        watermark[225] <= 18'b111111111111111111;
        watermark[226] <= 18'b111111111111111111;
        watermark[227] <= 18'b111111111111111111;
        watermark[228] <= 18'b111111111111111111;
        watermark[229] <= 18'b111111111111111111;
        watermark[230] <= 18'b111111111111111111;
        watermark[231] <= 18'b111111111111111111;
        watermark[232] <= 18'b111111111111111111;
        watermark[233] <= 18'b111111111111111111;
        watermark[234] <= 18'b111111111111111111;
        watermark[235] <= 18'b111111111111111111;
        watermark[236] <= 18'b111111111111111111;
        watermark[237] <= 18'b111111111111111111;
        watermark[238] <= 18'b111111111111111111;
        watermark[239] <= 18'b111111111111111111;
        watermark[240] <= 18'b111111111111111111;
        watermark[241] <= 18'b111111111111111111;
        watermark[242] <= 18'b111111111111111111;
        watermark[243] <= 18'b111111111111111111;
        watermark[244] <= 18'b111111111111111111;
        watermark[245] <= 18'b111111111111111111;
        watermark[246] <= 18'b111111111111111111;
        watermark[247] <= 18'b111111111111111111;
        watermark[248] <= 18'b111111111111111111;
        watermark[249] <= 18'b111111111111111111;
        watermark[250] <= 18'b111111111111111111;
        watermark[251] <= 18'b111111111111111111;
        watermark[252] <= 18'b111111111111111111;
        watermark[253] <= 18'b111111111111111111;
        watermark[254] <= 18'b111111111111111111;
        watermark[255] <= 18'b111111111111111111;
        watermark[256] <= 18'b111111111111111111;
        watermark[257] <= 18'b111111111111111111;
        watermark[258] <= 18'b111111111111111111;
        watermark[259] <= 18'b111111111111111111;
        watermark[260] <= 18'b111111111111111111;
        watermark[261] <= 18'b111111111111111111;
        watermark[262] <= 18'b111111111111111111;
        watermark[263] <= 18'b111111111111111111;
        watermark[264] <= 18'b111111111111111111;
        watermark[265] <= 18'b111111111111111111;
        watermark[266] <= 18'b111111111111111111;
        watermark[267] <= 18'b111111111111111111;
        watermark[268] <= 18'b111111111111111111;
        watermark[269] <= 18'b111111111111111111;
        watermark[270] <= 18'b111111111111111111;
        watermark[271] <= 18'b111111111111111111;
        watermark[272] <= 18'b111111111111111111;
        watermark[273] <= 18'b111111111111111111;
        watermark[274] <= 18'b111111111111111111;
        watermark[275] <= 18'b111111111111111111;
        watermark[276] <= 18'b111111111111111111;
        watermark[277] <= 18'b111111111111111111;
        watermark[278] <= 18'b111111111111111111;
        watermark[279] <= 18'b111111111111111111;
        watermark[280] <= 18'b111111111111111111;
        watermark[281] <= 18'b111111111111111111;
        watermark[282] <= 18'b111111111111111111;
        watermark[283] <= 18'b111111111111111111;
        watermark[284] <= 18'b111111111111111111;
        watermark[285] <= 18'b111111111111111111;
        watermark[286] <= 18'b111111111111111111;
        watermark[287] <= 18'b111111111111111111;
        watermark[288] <= 18'b111111111111111111;
        watermark[289] <= 18'b111111111111111111;
        watermark[290] <= 18'b111111111111111111;
        watermark[291] <= 18'b111111111111111111;
        watermark[292] <= 18'b111111111111111111;
        watermark[293] <= 18'b111111111111111111;
        watermark[294] <= 18'b111111111111111111;
        watermark[295] <= 18'b111111111111111111;
        watermark[296] <= 18'b111111111111111111;
        watermark[297] <= 18'b111111111111111111;
        watermark[298] <= 18'b111111111111111111;
        watermark[299] <= 18'b111111111111111111;
        watermark[300] <= 18'b111111111111111111;
        watermark[301] <= 18'b111111111111111111;
        watermark[302] <= 18'b111111111111111111;
        watermark[303] <= 18'b111111111111111111;
        watermark[304] <= 18'b111111111111110000;
        watermark[305] <= 18'b111111111111111111;
        watermark[306] <= 18'b110000111111111111;
        watermark[307] <= 18'b111111111111111111;
        watermark[308] <= 18'b111111111111111111;
        watermark[309] <= 18'b111111111111111111;
        watermark[310] <= 18'b111111111111111111;
        watermark[311] <= 18'b111111111111111111;
        watermark[312] <= 18'b111111111111111111;
        watermark[313] <= 18'b111111111111111111;
        watermark[314] <= 18'b111111111111111111;
        watermark[315] <= 18'b111111111110000000;
        watermark[316] <= 18'b001111111111111111;
        watermark[317] <= 18'b111100000000111111;
        watermark[318] <= 18'b111111111111111111;
        watermark[319] <= 18'b111111111111111111;
        watermark[320] <= 18'b111111111111111111;
        watermark[321] <= 18'b111111111111111111;
        watermark[322] <= 18'b111111111111111111;
        watermark[323] <= 18'b111111111111111111;
        watermark[324] <= 18'b111111111111111111;
        watermark[325] <= 18'b111111111111111111;
        watermark[326] <= 18'b111111111110000000;
        watermark[327] <= 18'b000001111111111111;
        watermark[328] <= 18'b111110000000000001;
        watermark[329] <= 18'b111111111111111111;
        watermark[330] <= 18'b111111111111111111;
        watermark[331] <= 18'b111111111111111111;
        watermark[332] <= 18'b111111111111111111;
        watermark[333] <= 18'b111111111111111111;
        watermark[334] <= 18'b111111111111111111;
        watermark[335] <= 18'b111111111111111111;
        watermark[336] <= 18'b111111111111111111;
        watermark[337] <= 18'b111111111110000000;
        watermark[338] <= 18'b000000011111111111;
        watermark[339] <= 18'b111111100000000000;
        watermark[340] <= 18'b000111111111111111;
        watermark[341] <= 18'b111111111111111111;
        watermark[342] <= 18'b111111111111111111;
        watermark[343] <= 18'b111111111111111111;
        watermark[344] <= 18'b111111111111111111;
        watermark[345] <= 18'b111111111111111111;
        watermark[346] <= 18'b111111111111111111;
        watermark[347] <= 18'b111111111111111111;
        watermark[348] <= 18'b111111111110000000;
        watermark[349] <= 18'b000000000011111111;
        watermark[350] <= 18'b111111110000000000;
        watermark[351] <= 18'b000000011111111111;
        watermark[352] <= 18'b111111111111111111;
        watermark[353] <= 18'b111111111111111111;
        watermark[354] <= 18'b111111111111111111;
        watermark[355] <= 18'b111111111111111111;
        watermark[356] <= 18'b111111111111111111;
        watermark[357] <= 18'b111111111111111111;
        watermark[358] <= 18'b111111111111111111;
        watermark[359] <= 18'b111111111111000000;
        watermark[360] <= 18'b000000000000111111;
        watermark[361] <= 18'b111111111100000000;
        watermark[362] <= 18'b000000000011111111;
        watermark[363] <= 18'b111111111111111111;
        watermark[364] <= 18'b111111111111111111;
        watermark[365] <= 18'b111111111111111111;
        watermark[366] <= 18'b111111111111111111;
        watermark[367] <= 18'b111111111111111111;
        watermark[368] <= 18'b111111111111111111;
        watermark[369] <= 18'b111111111111111111;
        watermark[370] <= 18'b111111111111100000;
        watermark[371] <= 18'b000000000000001111;
        watermark[372] <= 18'b111111111110000000;
        watermark[373] <= 18'b000000000000011111;
        watermark[374] <= 18'b111111111111111111;
        watermark[375] <= 18'b111111111111111111;
        watermark[376] <= 18'b111111111111111111;
        watermark[377] <= 18'b111111111111111111;
        watermark[378] <= 18'b111111111111111111;
        watermark[379] <= 18'b111111111111111111;
        watermark[380] <= 18'b111111111111111111;
        watermark[381] <= 18'b111111111111110000;
        watermark[382] <= 18'b000000000000000001;
        watermark[383] <= 18'b111111111111100000;
        watermark[384] <= 18'b000000000000000011;
        watermark[385] <= 18'b111111111111111111;
        watermark[386] <= 18'b111111111111111111;
        watermark[387] <= 18'b111111111111111111;
        watermark[388] <= 18'b111111111111111111;
        watermark[389] <= 18'b111111111111111111;
        watermark[390] <= 18'b111111111111111111;
        watermark[391] <= 18'b111111111111111111;
        watermark[392] <= 18'b111111111111111000;
        watermark[393] <= 18'b000000000000000000;
        watermark[394] <= 18'b011111111111111000;
        watermark[395] <= 18'b000000000000000000;
        watermark[396] <= 18'b011111111111111111;
        watermark[397] <= 18'b111111111111111111;
        watermark[398] <= 18'b111111111111111111;
        watermark[399] <= 18'b111111111111111111;
        watermark[400] <= 18'b111111111111111111;
        watermark[401] <= 18'b111111111111111111;
        watermark[402] <= 18'b111111111111111111;
        watermark[403] <= 18'b111111111111111100;
        watermark[404] <= 18'b000000000000000000;
        watermark[405] <= 18'b000111111111111110;
        watermark[406] <= 18'b000000000000000000;
        watermark[407] <= 18'b000011111111111111;
        watermark[408] <= 18'b111111111111111111;
        watermark[409] <= 18'b111111111111111111;
        watermark[410] <= 18'b111111111111111111;
        watermark[411] <= 18'b111111111111111111;
        watermark[412] <= 18'b111111111111111111;
        watermark[413] <= 18'b111111111111111111;
        watermark[414] <= 18'b111111111111111111;
        watermark[415] <= 18'b000000000000000000;
        watermark[416] <= 18'b000000111111111111;
        watermark[417] <= 18'b000000000000000000;
        watermark[418] <= 18'b000000111111111111;
        watermark[419] <= 18'b111111111111111111;
        watermark[420] <= 18'b111111111111111111;
        watermark[421] <= 18'b111111111111111111;
        watermark[422] <= 18'b111111111111111111;
        watermark[423] <= 18'b111111111111111111;
        watermark[424] <= 18'b111111111111111111;
        watermark[425] <= 18'b111111111111111111;
        watermark[426] <= 18'b100000000000000000;
        watermark[427] <= 18'b000000001111111111;
        watermark[428] <= 18'b110000000000000000;
        watermark[429] <= 18'b000000000111111111;
        watermark[430] <= 18'b111111111111111111;
        watermark[431] <= 18'b111111111111111111;
        watermark[432] <= 18'b111111111111111111;
        watermark[433] <= 18'b111111111111111111;
        watermark[434] <= 18'b111111111111111111;
        watermark[435] <= 18'b111111111111111111;
        watermark[436] <= 18'b111111111111111111;
        watermark[437] <= 18'b110000000000000000;
        watermark[438] <= 18'b000000000011111111;
        watermark[439] <= 18'b111100000000000000;
        watermark[440] <= 18'b000000000000111111;
        watermark[441] <= 18'b111111111111111111;
        watermark[442] <= 18'b111111111111111111;
        watermark[443] <= 18'b111111111111111111;
        watermark[444] <= 18'b111111111111111111;
        watermark[445] <= 18'b111111111111111111;
        watermark[446] <= 18'b111111111111111111;
        watermark[447] <= 18'b111111111111111111;
        watermark[448] <= 18'b111100000000000000;
        watermark[449] <= 18'b000000000000111111;
        watermark[450] <= 18'b111110000000000000;
        watermark[451] <= 18'b000000000000001111;
        watermark[452] <= 18'b111111111111111111;
        watermark[453] <= 18'b111111111111111111;
        watermark[454] <= 18'b111111111111111111;
        watermark[455] <= 18'b111111111111111111;
        watermark[456] <= 18'b111111111111111111;
        watermark[457] <= 18'b111111111111111111;
        watermark[458] <= 18'b111111111111111111;
        watermark[459] <= 18'b111111000000000000;
        watermark[460] <= 18'b000000000000000111;
        watermark[461] <= 18'b111111100000000000;
        watermark[462] <= 18'b000000000000000011;
        watermark[463] <= 18'b111111111111111111;
        watermark[464] <= 18'b111111111111111111;
        watermark[465] <= 18'b111111111111111111;
        watermark[466] <= 18'b111111111111111111;
        watermark[467] <= 18'b111111111111111111;
        watermark[468] <= 18'b111111111111111111;
        watermark[469] <= 18'b111111111111111111;
        watermark[470] <= 18'b111111100000000000;
        watermark[471] <= 18'b000000000000000001;
        watermark[472] <= 18'b111111111000000000;
        watermark[473] <= 18'b000000000000000000;
        watermark[474] <= 18'b011111111111111111;
        watermark[475] <= 18'b111111111111111111;
        watermark[476] <= 18'b111111111111111111;
        watermark[477] <= 18'b111111111111111111;
        watermark[478] <= 18'b111111111111111111;
        watermark[479] <= 18'b111111111111111111;
        watermark[480] <= 18'b111111111111111111;
        watermark[481] <= 18'b111111111000000000;
        watermark[482] <= 18'b000000000000000000;
        watermark[483] <= 18'b011111111110000000;
        watermark[484] <= 18'b000000000000000000;
        watermark[485] <= 18'b000111111111111111;
        watermark[486] <= 18'b111111111111111111;
        watermark[487] <= 18'b111111111111111111;
        watermark[488] <= 18'b111111111111111111;
        watermark[489] <= 18'b111111111111111111;
        watermark[490] <= 18'b111111111111111111;
        watermark[491] <= 18'b111111111111111111;
        watermark[492] <= 18'b111111111110000000;
        watermark[493] <= 18'b000000000000000000;
        watermark[494] <= 18'b000111111111100000;
        watermark[495] <= 18'b000000000000000000;
        watermark[496] <= 18'b000001111111111111;
        watermark[497] <= 18'b111111111111111111;
        watermark[498] <= 18'b111111111111111111;
        watermark[499] <= 18'b111111111111111111;
        watermark[500] <= 18'b111111111111111111;
        watermark[501] <= 18'b111111111111111111;
        watermark[502] <= 18'b111111111111111111;
        watermark[503] <= 18'b111111111111100000;
        watermark[504] <= 18'b000000000000000000;
        watermark[505] <= 18'b000000111111110000;
        watermark[506] <= 18'b000000000000000000;
        watermark[507] <= 18'b000000011111111111;
        watermark[508] <= 18'b111111111111111111;
        watermark[509] <= 18'b111111111111111111;
        watermark[510] <= 18'b111111111111111111;
        watermark[511] <= 18'b111111111111111111;
        watermark[512] <= 18'b111111111111111111;
        watermark[513] <= 18'b111111111111111111;
        watermark[514] <= 18'b111111111111111000;
        watermark[515] <= 18'b000000000000000000;
        watermark[516] <= 18'b000000001111111100;
        watermark[517] <= 18'b000000000000000000;
        watermark[518] <= 18'b000000000111111111;
        watermark[519] <= 18'b111111111111111111;
        watermark[520] <= 18'b111111111111111111;
        watermark[521] <= 18'b111111111111111111;
        watermark[522] <= 18'b111111111111111111;
        watermark[523] <= 18'b111111111111111111;
        watermark[524] <= 18'b111111111111111100;
        watermark[525] <= 18'b111111111111111100;
        watermark[526] <= 18'b000000000000000000;
        watermark[527] <= 18'b000000000011111111;
        watermark[528] <= 18'b000000000000000000;
        watermark[529] <= 18'b000000000001111111;
        watermark[530] <= 18'b111111111100111111;
        watermark[531] <= 18'b111111111111111111;
        watermark[532] <= 18'b111111111111111111;
        watermark[533] <= 18'b111111111111111111;
        watermark[534] <= 18'b111111111111111111;
        watermark[535] <= 18'b111111111111111110;
        watermark[536] <= 18'b000111111111111111;
        watermark[537] <= 18'b000000000000000000;
        watermark[538] <= 18'b000000000000111111;
        watermark[539] <= 18'b110000000000000000;
        watermark[540] <= 18'b000000000000011111;
        watermark[541] <= 18'b111111111110000111;
        watermark[542] <= 18'b111111111111111111;
        watermark[543] <= 18'b111111111111111111;
        watermark[544] <= 18'b111111111111111111;
        watermark[545] <= 18'b111111111111111111;
        watermark[546] <= 18'b111111111111111111;
        watermark[547] <= 18'b000000111111111111;
        watermark[548] <= 18'b110000000000000000;
        watermark[549] <= 18'b000000000000001111;
        watermark[550] <= 18'b111100000000000000;
        watermark[551] <= 18'b000000000000000111;
        watermark[552] <= 18'b111111111111000000;
        watermark[553] <= 18'b111111111111111111;
        watermark[554] <= 18'b111111111111111111;
        watermark[555] <= 18'b111111111111111111;
        watermark[556] <= 18'b111111111111111111;
        watermark[557] <= 18'b111111111111111111;
        watermark[558] <= 18'b110000000111111111;
        watermark[559] <= 18'b111100000000000000;
        watermark[560] <= 18'b000000000000000011;
        watermark[561] <= 18'b111111000000000000;
        watermark[562] <= 18'b000000000000000001;
        watermark[563] <= 18'b111111111111100000;
        watermark[564] <= 18'b001111111111111111;
        watermark[565] <= 18'b111111111111111111;
        watermark[566] <= 18'b111111111111111111;
        watermark[567] <= 18'b111111111111111111;
        watermark[568] <= 18'b111111111111111111;
        watermark[569] <= 18'b111000000001111111;
        watermark[570] <= 18'b111111100000000000;
        watermark[571] <= 18'b000000000000000000;
        watermark[572] <= 18'b111111100000000000;
        watermark[573] <= 18'b000000000000000000;
        watermark[574] <= 18'b011111111111110000;
        watermark[575] <= 18'b000001111111111111;
        watermark[576] <= 18'b111111111111111111;
        watermark[577] <= 18'b111111111111111111;
        watermark[578] <= 18'b111111111111111111;
        watermark[579] <= 18'b111111111111111111;
        watermark[580] <= 18'b111100000000001111;
        watermark[581] <= 18'b111111111000000000;
        watermark[582] <= 18'b000000000000000000;
        watermark[583] <= 18'b000111111000000000;
        watermark[584] <= 18'b000000000000000000;
        watermark[585] <= 18'b000111111111111100;
        watermark[586] <= 18'b000000001111111111;
        watermark[587] <= 18'b111111111111111111;
        watermark[588] <= 18'b111111111111111111;
        watermark[589] <= 18'b111111111111111111;
        watermark[590] <= 18'b111111111111111111;
        watermark[591] <= 18'b111110000000000001;
        watermark[592] <= 18'b111111111110000000;
        watermark[593] <= 18'b000000000000000000;
        watermark[594] <= 18'b000001111110000000;
        watermark[595] <= 18'b000000000000000000;
        watermark[596] <= 18'b000001111111111110;
        watermark[597] <= 18'b000000000001111111;
        watermark[598] <= 18'b111111111111111111;
        watermark[599] <= 18'b111111111111111111;
        watermark[600] <= 18'b111111111111111111;
        watermark[601] <= 18'b111111111111111111;
        watermark[602] <= 18'b111111100000000000;
        watermark[603] <= 18'b001111111111100000;
        watermark[604] <= 18'b000000000000000000;
        watermark[605] <= 18'b000000011111100000;
        watermark[606] <= 18'b000000000000000000;
        watermark[607] <= 18'b000000011111111111;
        watermark[608] <= 18'b000000000000011111;
        watermark[609] <= 18'b111111111111111111;
        watermark[610] <= 18'b111111111111111111;
        watermark[611] <= 18'b111111111111111111;
        watermark[612] <= 18'b111111111111111111;
        watermark[613] <= 18'b111111110000000000;
        watermark[614] <= 18'b000011111111111000;
        watermark[615] <= 18'b000000000000000000;
        watermark[616] <= 18'b000000000111111000;
        watermark[617] <= 18'b000000000000000000;
        watermark[618] <= 18'b000000000111111111;
        watermark[619] <= 18'b110000000000000011;
        watermark[620] <= 18'b111111111111111111;
        watermark[621] <= 18'b111111111111111111;
        watermark[622] <= 18'b111111111111111111;
        watermark[623] <= 18'b111111111111111111;
        watermark[624] <= 18'b111111111000000000;
        watermark[625] <= 18'b000000011111111110;
        watermark[626] <= 18'b000000000000000000;
        watermark[627] <= 18'b000000000001111110;
        watermark[628] <= 18'b000000000000000000;
        watermark[629] <= 18'b000000000001111111;
        watermark[630] <= 18'b111000000000000000;
        watermark[631] <= 18'b011111111111111111;
        watermark[632] <= 18'b111111111111111111;
        watermark[633] <= 18'b111111111111111111;
        watermark[634] <= 18'b111111111111111111;
        watermark[635] <= 18'b111111111110000000;
        watermark[636] <= 18'b000000000011111111;
        watermark[637] <= 18'b110000000000000000;
        watermark[638] <= 18'b000000000000011111;
        watermark[639] <= 18'b100000000000000000;
        watermark[640] <= 18'b000000000000111111;
        watermark[641] <= 18'b111100000000000000;
        watermark[642] <= 18'b000111111111111111;
        watermark[643] <= 18'b111111111111111111;
        watermark[644] <= 18'b111111111111111111;
        watermark[645] <= 18'b111111111111111111;
        watermark[646] <= 18'b111111111111000000;
        watermark[647] <= 18'b000000000000011111;
        watermark[648] <= 18'b111100000000000000;
        watermark[649] <= 18'b000000000000000111;
        watermark[650] <= 18'b111000000000000000;
        watermark[651] <= 18'b000000000000001111;
        watermark[652] <= 18'b111110000000000000;
        watermark[653] <= 18'b000000111111111111;
        watermark[654] <= 18'b111111111111111111;
        watermark[655] <= 18'b111111111111111111;
        watermark[656] <= 18'b111111111111111111;
        watermark[657] <= 18'b111111111111110000;
        watermark[658] <= 18'b000000000000000111;
        watermark[659] <= 18'b111111000000000000;
        watermark[660] <= 18'b000000000000000001;
        watermark[661] <= 18'b111110000000000000;
        watermark[662] <= 18'b000000000000000011;
        watermark[663] <= 18'b111111100000000000;
        watermark[664] <= 18'b000000001111111111;
        watermark[665] <= 18'b111111111111111111;
        watermark[666] <= 18'b111111111111111111;
        watermark[667] <= 18'b111111111111111111;
        watermark[668] <= 18'b111111111111111000;
        watermark[669] <= 18'b000000000000000000;
        watermark[670] <= 18'b111111111000000000;
        watermark[671] <= 18'b000000000000000000;
        watermark[672] <= 18'b011111100000000000;
        watermark[673] <= 18'b000000000000000001;
        watermark[674] <= 18'b111111110000000000;
        watermark[675] <= 18'b000000000001111111;
        watermark[676] <= 18'b111111111111111111;
        watermark[677] <= 18'b111111111111111111;
        watermark[678] <= 18'b111111111111111111;
        watermark[679] <= 18'b111111111111111110;
        watermark[680] <= 18'b000000000000000000;
        watermark[681] <= 18'b000111111110000000;
        watermark[682] <= 18'b000000000000000000;
        watermark[683] <= 18'b000111110000000000;
        watermark[684] <= 18'b000000000000000000;
        watermark[685] <= 18'b011111111000000000;
        watermark[686] <= 18'b000000000000011111;
        watermark[687] <= 18'b111111111111111111;
        watermark[688] <= 18'b111111111111111111;
        watermark[689] <= 18'b111111111111111111;
        watermark[690] <= 18'b111111111111111111;
        watermark[691] <= 18'b100000000000000000;
        watermark[692] <= 18'b000001111111100000;
        watermark[693] <= 18'b000000000000000000;
        watermark[694] <= 18'b000000111100000000;
        watermark[695] <= 18'b000000000000000000;
        watermark[696] <= 18'b000111111110000000;
        watermark[697] <= 18'b000000000000000111;
        watermark[698] <= 18'b111111111111111111;
        watermark[699] <= 18'b111111111111111111;
        watermark[700] <= 18'b111111111111111111;
        watermark[701] <= 18'b111111111111111111;
        watermark[702] <= 18'b110000000000000000;
        watermark[703] <= 18'b000000001111111100;
        watermark[704] <= 18'b000000000000000000;
        watermark[705] <= 18'b000000001111000000;
        watermark[706] <= 18'b000000000000000000;
        watermark[707] <= 18'b000011111111000000;
        watermark[708] <= 18'b000000000000000000;
        watermark[709] <= 18'b111111111111111111;
        watermark[710] <= 18'b111111111111111111;
        watermark[711] <= 18'b111111111111111111;
        watermark[712] <= 18'b111111111111111111;
        watermark[713] <= 18'b111100000000000000;
        watermark[714] <= 18'b000000000001111111;
        watermark[715] <= 18'b000000000000000000;
        watermark[716] <= 18'b000000000011110000;
        watermark[717] <= 18'b000000000000000000;
        watermark[718] <= 18'b000000111111100000;
        watermark[719] <= 18'b000000000000000000;
        watermark[720] <= 18'b001111111111111111;
        watermark[721] <= 18'b111111111111111111;
        watermark[722] <= 18'b111111111111111111;
        watermark[723] <= 18'b111111111111111111;
        watermark[724] <= 18'b111111000000000000;
        watermark[725] <= 18'b000000000000011111;
        watermark[726] <= 18'b110000000000000000;
        watermark[727] <= 18'b000000000000111100;
        watermark[728] <= 18'b000000000000000000;
        watermark[729] <= 18'b000000001111110000;
        watermark[730] <= 18'b000000000000000000;
        watermark[731] <= 18'b000011111111111111;
        watermark[732] <= 18'b111111111111111111;
        watermark[733] <= 18'b111111111111111111;
        watermark[734] <= 18'b111111111111111111;
        watermark[735] <= 18'b111111110000000000;
        watermark[736] <= 18'b000000000000000011;
        watermark[737] <= 18'b111110000000000000;
        watermark[738] <= 18'b000000000000001111;
        watermark[739] <= 18'b000000000000000000;
        watermark[740] <= 18'b000000000111111100;
        watermark[741] <= 18'b000000000000000000;
        watermark[742] <= 18'b000000111111111111;
        watermark[743] <= 18'b111111111111111111;
        watermark[744] <= 18'b111111111111111111;
        watermark[745] <= 18'b111111111111111111;
        watermark[746] <= 18'b111111111100000000;
        watermark[747] <= 18'b000000000000000000;
        watermark[748] <= 18'b011111100000000000;
        watermark[749] <= 18'b000000000000000011;
        watermark[750] <= 18'b110000000000000000;
        watermark[751] <= 18'b000000000001111110;
        watermark[752] <= 18'b000000000000000000;
        watermark[753] <= 18'b000000001111111111;
        watermark[754] <= 18'b111111111111111111;
        watermark[755] <= 18'b111111111111111111;
        watermark[756] <= 18'b111111111111111111;
        watermark[757] <= 18'b111111111110000000;
        watermark[758] <= 18'b000000000000000000;
        watermark[759] <= 18'b000111111100000000;
        watermark[760] <= 18'b000000000000000000;
        watermark[761] <= 18'b111100000000000000;
        watermark[762] <= 18'b000000000000111111;
        watermark[763] <= 18'b000000000000000000;
        watermark[764] <= 18'b000000000011111111;
        watermark[765] <= 18'b111111111111111111;
        watermark[766] <= 18'b111111111111111111;
        watermark[767] <= 18'b111111111111111111;
        watermark[768] <= 18'b111111111111100000;
        watermark[769] <= 18'b000000000000000000;
        watermark[770] <= 18'b000000111111000000;
        watermark[771] <= 18'b000000000000000000;
        watermark[772] <= 18'b001111000000000000;
        watermark[773] <= 18'b000000000000001111;
        watermark[774] <= 18'b110000000000000000;
        watermark[775] <= 18'b000000000000111111;
        watermark[776] <= 18'b111111111111111111;
        watermark[777] <= 18'b111111111111111111;
        watermark[778] <= 18'b111111111111111111;
        watermark[779] <= 18'b111111111111111000;
        watermark[780] <= 18'b000000000000000000;
        watermark[781] <= 18'b000000000111110000;
        watermark[782] <= 18'b000000000000000000;
        watermark[783] <= 18'b000011110000000000;
        watermark[784] <= 18'b000000000000000111;
        watermark[785] <= 18'b111000000000000000;
        watermark[786] <= 18'b000000000000001111;
        watermark[787] <= 18'b111111111111111111;
        watermark[788] <= 18'b111111111111111111;
        watermark[789] <= 18'b111111111111111111;
        watermark[790] <= 18'b111111111111111111;
        watermark[791] <= 18'b000000000000000000;
        watermark[792] <= 18'b000000000001111110;
        watermark[793] <= 18'b000000000000000000;
        watermark[794] <= 18'b000000111100000000;
        watermark[795] <= 18'b000000000000000001;
        watermark[796] <= 18'b111100000000000000;
        watermark[797] <= 18'b000000000000000011;
        watermark[798] <= 18'b111111111111111111;
        watermark[799] <= 18'b111111111111111111;
        watermark[800] <= 18'b111111111111111111;
        watermark[801] <= 18'b111111111111111111;
        watermark[802] <= 18'b110000000000000000;
        watermark[803] <= 18'b000000000000001111;
        watermark[804] <= 18'b100000000000000000;
        watermark[805] <= 18'b000000001111000000;
        watermark[806] <= 18'b000000000000000000;
        watermark[807] <= 18'b011111000000000000;
        watermark[808] <= 18'b000000000000000000;
        watermark[809] <= 18'b111111111111111111;
        watermark[810] <= 18'b111111111111111111;
        watermark[811] <= 18'b111111111111111111;
        watermark[812] <= 18'b111111111111111111;
        watermark[813] <= 18'b111100000000000000;
        watermark[814] <= 18'b000000000000000001;
        watermark[815] <= 18'b111100000000000000;
        watermark[816] <= 18'b000000000011110000;
        watermark[817] <= 18'b000000000000000000;
        watermark[818] <= 18'b001111100000000000;
        watermark[819] <= 18'b000000000000000000;
        watermark[820] <= 18'b001111111111111111;
        watermark[821] <= 18'b111111111111111111;
        watermark[822] <= 18'b111111111111111111;
        watermark[823] <= 18'b111111111111111111;
        watermark[824] <= 18'b111111000000000000;
        watermark[825] <= 18'b000000000000000000;
        watermark[826] <= 18'b011111000000000000;
        watermark[827] <= 18'b000000000000111100;
        watermark[828] <= 18'b000000000000000000;
        watermark[829] <= 18'b000011111000000000;
        watermark[830] <= 18'b000000000000000000;
        watermark[831] <= 18'b000011111111111111;
        watermark[832] <= 18'b111111111111111111;
        watermark[833] <= 18'b111111111111111111;
        watermark[834] <= 18'b111111111111111111;
        watermark[835] <= 18'b111111110000000000;
        watermark[836] <= 18'b000000000000000000;
        watermark[837] <= 18'b000011111000000000;
        watermark[838] <= 18'b000000000000001111;
        watermark[839] <= 18'b000000000000000000;
        watermark[840] <= 18'b000001111100000000;
        watermark[841] <= 18'b000000000000000000;
        watermark[842] <= 18'b000000111111111111;
        watermark[843] <= 18'b111111111111111111;
        watermark[844] <= 18'b111111111111111111;
        watermark[845] <= 18'b111111111111111111;
        watermark[846] <= 18'b111111111110000000;
        watermark[847] <= 18'b000000000000000000;
        watermark[848] <= 18'b000000011110000000;
        watermark[849] <= 18'b000000000000000011;
        watermark[850] <= 18'b110000000000000000;
        watermark[851] <= 18'b000000011110000000;
        watermark[852] <= 18'b000000000000000000;
        watermark[853] <= 18'b000000011111111111;
        watermark[854] <= 18'b111111111111111111;
        watermark[855] <= 18'b111111111111111111;
        watermark[856] <= 18'b111111111111111111;
        watermark[857] <= 18'b111111111111100000;
        watermark[858] <= 18'b000000000000000000;
        watermark[859] <= 18'b000000000111110000;
        watermark[860] <= 18'b000000000000000000;
        watermark[861] <= 18'b111100000000000000;
        watermark[862] <= 18'b000000001111100000;
        watermark[863] <= 18'b000000000000000000;
        watermark[864] <= 18'b000000000111111111;
        watermark[865] <= 18'b111111111111111111;
        watermark[866] <= 18'b111111111111111111;
        watermark[867] <= 18'b111111111111111111;
        watermark[868] <= 18'b111111111111111100;
        watermark[869] <= 18'b000000000000000000;
        watermark[870] <= 18'b000000000000111100;
        watermark[871] <= 18'b000000000000000000;
        watermark[872] <= 18'b001111000000000000;
        watermark[873] <= 18'b000000000011110000;
        watermark[874] <= 18'b000000000000000000;
        watermark[875] <= 18'b000000000011111111;
        watermark[876] <= 18'b111111111111111111;
        watermark[877] <= 18'b111111111111111111;
        watermark[878] <= 18'b111111111111111111;
        watermark[879] <= 18'b111111111111111111;
        watermark[880] <= 18'b000000000000000000;
        watermark[881] <= 18'b000000000000000111;
        watermark[882] <= 18'b100000000000000000;
        watermark[883] <= 18'b000011110000000000;
        watermark[884] <= 18'b000000000001111000;
        watermark[885] <= 18'b000000000000000000;
        watermark[886] <= 18'b000000000000111111;
        watermark[887] <= 18'b111111111111111111;
        watermark[888] <= 18'b111111111111111111;
        watermark[889] <= 18'b111111111111111111;
        watermark[890] <= 18'b111111111111111111;
        watermark[891] <= 18'b111000000000000000;
        watermark[892] <= 18'b000000000000000001;
        watermark[893] <= 18'b111000000000000000;
        watermark[894] <= 18'b000000111100000000;
        watermark[895] <= 18'b000000000000111110;
        watermark[896] <= 18'b000000000000000000;
        watermark[897] <= 18'b000000000000011111;
        watermark[898] <= 18'b111111111111111111;
        watermark[899] <= 18'b111111111111111111;
        watermark[900] <= 18'b111111111111111111;
        watermark[901] <= 18'b111111111111111111;
        watermark[902] <= 18'b111110000000000000;
        watermark[903] <= 18'b000000000000000000;
        watermark[904] <= 18'b001111000000000000;
        watermark[905] <= 18'b000000001111000000;
        watermark[906] <= 18'b000000000000001111;
        watermark[907] <= 18'b000000000000000000;
        watermark[908] <= 18'b000000000000001111;
        watermark[909] <= 18'b111111111111111111;
        watermark[910] <= 18'b111111111111111111;
        watermark[911] <= 18'b111111111111111111;
        watermark[912] <= 18'b111111111111111111;
        watermark[913] <= 18'b111111110000000000;
        watermark[914] <= 18'b000000000000000000;
        watermark[915] <= 18'b000011111000000000;
        watermark[916] <= 18'b000000000011110000;
        watermark[917] <= 18'b000000000000000111;
        watermark[918] <= 18'b110000000000000000;
        watermark[919] <= 18'b000000000000000011;
        watermark[920] <= 18'b111111111111111111;
        watermark[921] <= 18'b111111111111111111;
        watermark[922] <= 18'b111111111111111111;
        watermark[923] <= 18'b111111111111111111;
        watermark[924] <= 18'b111111111110000000;
        watermark[925] <= 18'b000000000000000000;
        watermark[926] <= 18'b000000011110000000;
        watermark[927] <= 18'b000000000000111100;
        watermark[928] <= 18'b000000000000000001;
        watermark[929] <= 18'b111000000000000000;
        watermark[930] <= 18'b000000000000000001;
        watermark[931] <= 18'b111111111111111111;
        watermark[932] <= 18'b111111111111111111;
        watermark[933] <= 18'b111111111111111111;
        watermark[934] <= 18'b111111111111111100;
        watermark[935] <= 18'b111111111111110000;
        watermark[936] <= 18'b000000000000000000;
        watermark[937] <= 18'b000000000011110000;
        watermark[938] <= 18'b000000000000001111;
        watermark[939] <= 18'b000000000000000000;
        watermark[940] <= 18'b111100000000000000;
        watermark[941] <= 18'b000000000000000000;
        watermark[942] <= 18'b111111111111110011;
        watermark[943] <= 18'b111111111111111111;
        watermark[944] <= 18'b111111111111111111;
        watermark[945] <= 18'b111111111111111111;
        watermark[946] <= 18'b000011111111111110;
        watermark[947] <= 18'b000000000000000000;
        watermark[948] <= 18'b000000000000111100;
        watermark[949] <= 18'b000000000000000011;
        watermark[950] <= 18'b110000000000000000;
        watermark[951] <= 18'b001111000000000000;
        watermark[952] <= 18'b000000000000000000;
        watermark[953] <= 18'b011111111111110000;
        watermark[954] <= 18'b111111111111111111;
        watermark[955] <= 18'b111111111111111111;
        watermark[956] <= 18'b111111111111111111;
        watermark[957] <= 18'b100000001111111111;
        watermark[958] <= 18'b110000000000000000;
        watermark[959] <= 18'b000000000000000111;
        watermark[960] <= 18'b100000000000000000;
        watermark[961] <= 18'b111100000000000000;
        watermark[962] <= 18'b000111100000000000;
        watermark[963] <= 18'b000000000000000000;
        watermark[964] <= 18'b001111111111110000;
        watermark[965] <= 18'b001111111111111111;
        watermark[966] <= 18'b111111111111111111;
        watermark[967] <= 18'b111111111111111111;
        watermark[968] <= 18'b111000000000111111;
        watermark[969] <= 18'b111110000000000000;
        watermark[970] <= 18'b000000000000000001;
        watermark[971] <= 18'b111000000000000000;
        watermark[972] <= 18'b001111000000000000;
        watermark[973] <= 18'b000011111000000000;
        watermark[974] <= 18'b000000000000000000;
        watermark[975] <= 18'b000111111111110000;
        watermark[976] <= 18'b000001111111111111;
        watermark[977] <= 18'b111111111111111111;
        watermark[978] <= 18'b111111111111111111;
        watermark[979] <= 18'b111110000000000111;
        watermark[980] <= 18'b111111111000000000;
        watermark[981] <= 18'b000000000000000000;
        watermark[982] <= 18'b001111000000000000;
        watermark[983] <= 18'b000011110000000000;
        watermark[984] <= 18'b000000111100000000;
        watermark[985] <= 18'b000000000000000000;
        watermark[986] <= 18'b000111111111110000;
        watermark[987] <= 18'b000000011111111111;
        watermark[988] <= 18'b111111111111111111;
        watermark[989] <= 18'b111111111111111111;
        watermark[990] <= 18'b111111100000000000;
        watermark[991] <= 18'b011111111111000000;
        watermark[992] <= 18'b000000000000000000;
        watermark[993] <= 18'b000011111000000000;
        watermark[994] <= 18'b000000111100000000;
        watermark[995] <= 18'b000000011111000000;
        watermark[996] <= 18'b000000000000000000;
        watermark[997] <= 18'b000011111111111000;
        watermark[998] <= 18'b000000000111111111;
        watermark[999] <= 18'b111111111111111111;
        watermark[1000] <= 18'b111111111111111111;
        watermark[1001] <= 18'b111111111000000000;
        watermark[1002] <= 18'b000001111111111000;
        watermark[1003] <= 18'b000000000000000000;
        watermark[1004] <= 18'b000000011110000000;
        watermark[1005] <= 18'b000000011111000000;
        watermark[1006] <= 18'b000000000111100000;
        watermark[1007] <= 18'b000000000000000000;
        watermark[1008] <= 18'b000001111111111000;
        watermark[1009] <= 18'b000000000001111111;
        watermark[1010] <= 18'b111111111111111111;
        watermark[1011] <= 18'b111111111111111111;
        watermark[1012] <= 18'b111111111110000000;
        watermark[1013] <= 18'b000000000111111111;
        watermark[1014] <= 18'b000000000000000000;
        watermark[1015] <= 18'b000000000011110000;
        watermark[1016] <= 18'b000000000111110000;
        watermark[1017] <= 18'b000000000011110000;
        watermark[1018] <= 18'b000000000000000000;
        watermark[1019] <= 18'b000001111111111000;
        watermark[1020] <= 18'b000000000000011111;
        watermark[1021] <= 18'b111111111111111111;
        watermark[1022] <= 18'b111111111111111111;
        watermark[1023] <= 18'b111111111111100000;
        watermark[1024] <= 18'b000000000000011111;
        watermark[1025] <= 18'b111100000000000000;
        watermark[1026] <= 18'b000000000000111100;
        watermark[1027] <= 18'b000000000001111110;
        watermark[1028] <= 18'b000000000000111100;
        watermark[1029] <= 18'b000000000000000000;
        watermark[1030] <= 18'b000000111111111000;
        watermark[1031] <= 18'b000000000000000111;
        watermark[1032] <= 18'b111111111111111111;
        watermark[1033] <= 18'b111111111111111111;
        watermark[1034] <= 18'b111111111111111000;
        watermark[1035] <= 18'b000000000000000011;
        watermark[1036] <= 18'b111111100000000000;
        watermark[1037] <= 18'b000000000000000111;
        watermark[1038] <= 18'b100000000000011111;
        watermark[1039] <= 18'b100000000000011110;
        watermark[1040] <= 18'b000000000000000000;
        watermark[1041] <= 18'b000000011111111000;
        watermark[1042] <= 18'b000000000000000001;
        watermark[1043] <= 18'b111111111111111111;
        watermark[1044] <= 18'b111111111111111111;
        watermark[1045] <= 18'b111111111111111110;
        watermark[1046] <= 18'b000000000000000000;
        watermark[1047] <= 18'b001111111110000000;
        watermark[1048] <= 18'b000000000000000001;
        watermark[1049] <= 18'b111100000000000111;
        watermark[1050] <= 18'b111000000000001111;
        watermark[1051] <= 18'b100000000000000000;
        watermark[1052] <= 18'b000000011111111100;
        watermark[1053] <= 18'b000000000000000000;
        watermark[1054] <= 18'b011111111111111111;
        watermark[1055] <= 18'b111111111111111111;
        watermark[1056] <= 18'b111111111111111111;
        watermark[1057] <= 18'b100000000000000000;
        watermark[1058] <= 18'b000000111111110000;
        watermark[1059] <= 18'b000000000000000000;
        watermark[1060] <= 18'b001111000000000001;
        watermark[1061] <= 18'b111110000000000011;
        watermark[1062] <= 18'b110000000000000000;
        watermark[1063] <= 18'b000000001111111100;
        watermark[1064] <= 18'b000000000000000000;
        watermark[1065] <= 18'b000111111111111111;
        watermark[1066] <= 18'b111111111111111111;
        watermark[1067] <= 18'b111111111111111111;
        watermark[1068] <= 18'b111000000000000000;
        watermark[1069] <= 18'b000000000011111111;
        watermark[1070] <= 18'b000000000000000000;
        watermark[1071] <= 18'b000011111000000000;
        watermark[1072] <= 18'b011111100000000001;
        watermark[1073] <= 18'b111100000000000000;
        watermark[1074] <= 18'b000000001111111100;
        watermark[1075] <= 18'b000000000000000000;
        watermark[1076] <= 18'b000001111111111111;
        watermark[1077] <= 18'b111111111111111111;
        watermark[1078] <= 18'b111111111111111111;
        watermark[1079] <= 18'b111111000000000000;
        watermark[1080] <= 18'b000000000000001111;
        watermark[1081] <= 18'b111000000000000000;
        watermark[1082] <= 18'b000000011111000000;
        watermark[1083] <= 18'b000111111000000000;
        watermark[1084] <= 18'b111110000000000000;
        watermark[1085] <= 18'b000000001111111100;
        watermark[1086] <= 18'b000000000000000000;
        watermark[1087] <= 18'b000000111111111111;
        watermark[1088] <= 18'b111111111111111111;
        watermark[1089] <= 18'b111111111111111111;
        watermark[1090] <= 18'b111111110000000000;
        watermark[1091] <= 18'b000000000000000001;
        watermark[1092] <= 18'b111111100000000000;
        watermark[1093] <= 18'b000000000111110000;
        watermark[1094] <= 18'b000001111110000000;
        watermark[1095] <= 18'b001111100000000000;
        watermark[1096] <= 18'b000000000111111110;
        watermark[1097] <= 18'b000000000000000000;
        watermark[1098] <= 18'b000000001111111111;
        watermark[1099] <= 18'b111111111111111111;
        watermark[1100] <= 18'b111111111111111111;
        watermark[1101] <= 18'b111111111100000000;
        watermark[1102] <= 18'b000000000000000000;
        watermark[1103] <= 18'b000111111110000000;
        watermark[1104] <= 18'b000000000000111110;
        watermark[1105] <= 18'b000000011111100000;
        watermark[1106] <= 18'b000111110000000000;
        watermark[1107] <= 18'b000000000111111110;
        watermark[1108] <= 18'b000000000000000000;
        watermark[1109] <= 18'b000000000011111111;
        watermark[1110] <= 18'b111111111111111111;
        watermark[1111] <= 18'b111111111111111111;
        watermark[1112] <= 18'b111111111111000000;
        watermark[1113] <= 18'b000000000000000000;
        watermark[1114] <= 18'b000000011111110000;
        watermark[1115] <= 18'b000000000000001111;
        watermark[1116] <= 18'b100000000111111000;
        watermark[1117] <= 18'b000011111100000000;
        watermark[1118] <= 18'b000000000011111110;
        watermark[1119] <= 18'b000000000000000000;
        watermark[1120] <= 18'b000000000000111111;
        watermark[1121] <= 18'b111111111111111111;
        watermark[1122] <= 18'b111111111111111111;
        watermark[1123] <= 18'b111111111111111000;
        watermark[1124] <= 18'b000000000000000000;
        watermark[1125] <= 18'b000000000001111111;
        watermark[1126] <= 18'b000000000000000001;
        watermark[1127] <= 18'b111100000001111110;
        watermark[1128] <= 18'b000000111110000000;
        watermark[1129] <= 18'b000000000011111110;
        watermark[1130] <= 18'b000000000000000000;
        watermark[1131] <= 18'b000000000000011111;
        watermark[1132] <= 18'b111111111111111111;
        watermark[1133] <= 18'b111111111111111111;
        watermark[1134] <= 18'b111111111111111110;
        watermark[1135] <= 18'b000000000000000000;
        watermark[1136] <= 18'b000000000000001111;
        watermark[1137] <= 18'b111100000000000000;
        watermark[1138] <= 18'b011111100000011111;
        watermark[1139] <= 18'b100000011111100000;
        watermark[1140] <= 18'b000000000011111111;
        watermark[1141] <= 18'b000000000000000000;
        watermark[1142] <= 18'b000000000000000111;
        watermark[1143] <= 18'b111111111111111111;
        watermark[1144] <= 18'b111111111111111111;
        watermark[1145] <= 18'b111111111111111111;
        watermark[1146] <= 18'b110000000000000000;
        watermark[1147] <= 18'b000000000000000000;
        watermark[1148] <= 18'b111111110000000000;
        watermark[1149] <= 18'b000011111000000111;
        watermark[1150] <= 18'b111000000111110000;
        watermark[1151] <= 18'b000000000011111111;
        watermark[1152] <= 18'b000000000000000000;
        watermark[1153] <= 18'b000000000000000011;
        watermark[1154] <= 18'b111111111111111111;
        watermark[1155] <= 18'b111111111111111111;
        watermark[1156] <= 18'b111111111111111111;
        watermark[1157] <= 18'b111100000000000000;
        watermark[1158] <= 18'b000000000000000000;
        watermark[1159] <= 18'b000011111110000000;
        watermark[1160] <= 18'b000000111111000001;
        watermark[1161] <= 18'b111110000011111100;
        watermark[1162] <= 18'b000000000001111111;
        watermark[1163] <= 18'b000000000000000000;
        watermark[1164] <= 18'b000000000000000000;
        watermark[1165] <= 18'b111111111111111111;
        watermark[1166] <= 18'b111111111111111111;
        watermark[1167] <= 18'b111111111111111111;
        watermark[1168] <= 18'b111111100000000000;
        watermark[1169] <= 18'b000000000000000000;
        watermark[1170] <= 18'b000000011111111000;
        watermark[1171] <= 18'b000000000111111000;
        watermark[1172] <= 18'b111111100001111110;
        watermark[1173] <= 18'b000000000001111111;
        watermark[1174] <= 18'b100000000000000000;
        watermark[1175] <= 18'b000000000000000000;
        watermark[1176] <= 18'b011111111111111111;
        watermark[1177] <= 18'b111111111111111111;
        watermark[1178] <= 18'b111111111111111111;
        watermark[1179] <= 18'b111111111000000000;
        watermark[1180] <= 18'b000000000000000000;
        watermark[1181] <= 18'b000000000001111111;
        watermark[1182] <= 18'b100000000001111110;
        watermark[1183] <= 18'b001111111100011111;
        watermark[1184] <= 18'b100000000001111111;
        watermark[1185] <= 18'b100000000000000000;
        watermark[1186] <= 18'b000000000000000000;
        watermark[1187] <= 18'b000111111111111111;
        watermark[1188] <= 18'b111111111111111111;
        watermark[1189] <= 18'b111111111111111111;
        watermark[1190] <= 18'b111111111111000000;
        watermark[1191] <= 18'b000000000000000000;
        watermark[1192] <= 18'b000000000000000111;
        watermark[1193] <= 18'b111110000000001111;
        watermark[1194] <= 18'b110011111111001111;
        watermark[1195] <= 18'b110000000001111111;
        watermark[1196] <= 18'b100000000000000000;
        watermark[1197] <= 18'b000000000000000000;
        watermark[1198] <= 18'b000011111111111111;
        watermark[1199] <= 18'b111111111111111111;
        watermark[1200] <= 18'b111111111111111111;
        watermark[1201] <= 18'b111111111111111000;
        watermark[1202] <= 18'b000000000000000000;
        watermark[1203] <= 18'b000000000000000000;
        watermark[1204] <= 18'b111111111000000011;
        watermark[1205] <= 18'b111110111111110111;
        watermark[1206] <= 18'b111100000001111111;
        watermark[1207] <= 18'b110000000000000000;
        watermark[1208] <= 18'b000000000000000000;
        watermark[1209] <= 18'b000001111111111111;
        watermark[1210] <= 18'b111111111111111111;
        watermark[1211] <= 18'b111111111111111111;
        watermark[1212] <= 18'b111111111111111111;
        watermark[1213] <= 18'b000000000000000000;
        watermark[1214] <= 18'b000000000000000000;
        watermark[1215] <= 18'b000011111111100000;
        watermark[1216] <= 18'b011111111111111111;
        watermark[1217] <= 18'b111110000001111111;
        watermark[1218] <= 18'b110000000000000000;
        watermark[1219] <= 18'b000000000000000000;
        watermark[1220] <= 18'b000000111111111111;
        watermark[1221] <= 18'b111111111111111111;
        watermark[1222] <= 18'b111111111111111111;
        watermark[1223] <= 18'b111111111111111111;
        watermark[1224] <= 18'b111000000000000000;
        watermark[1225] <= 18'b000000000000000000;
        watermark[1226] <= 18'b000000001111111110;
        watermark[1227] <= 18'b000111111111111111;
        watermark[1228] <= 18'b111111100001111111;
        watermark[1229] <= 18'b110000000000000000;
        watermark[1230] <= 18'b000000000000000000;
        watermark[1231] <= 18'b000000011111111111;
        watermark[1232] <= 18'b111111111111111111;
        watermark[1233] <= 18'b111111111111111111;
        watermark[1234] <= 18'b111111111111111111;
        watermark[1235] <= 18'b111111000000000000;
        watermark[1236] <= 18'b000000000000000000;
        watermark[1237] <= 18'b000000000001111111;
        watermark[1238] <= 18'b110000111111111111;
        watermark[1239] <= 18'b111111110001111111;
        watermark[1240] <= 18'b111000000000000000;
        watermark[1241] <= 18'b000000000000000000;
        watermark[1242] <= 18'b000000001111111111;
        watermark[1243] <= 18'b111111111111111111;
        watermark[1244] <= 18'b111111111111111111;
        watermark[1245] <= 18'b111111111111111111;
        watermark[1246] <= 18'b111111111000000000;
        watermark[1247] <= 18'b000000000000000000;
        watermark[1248] <= 18'b000000000000000111;
        watermark[1249] <= 18'b111111001111111111;
        watermark[1250] <= 18'b111111111101111111;
        watermark[1251] <= 18'b111000000000000000;
        watermark[1252] <= 18'b000000000000000000;
        watermark[1253] <= 18'b000000000111111111;
        watermark[1254] <= 18'b111111111111111111;
        watermark[1255] <= 18'b111111111111111111;
        watermark[1256] <= 18'b111111111111111111;
        watermark[1257] <= 18'b111111111111000000;
        watermark[1258] <= 18'b000000000000000000;
        watermark[1259] <= 18'b000000000000000000;
        watermark[1260] <= 18'b111111111111111111;
        watermark[1261] <= 18'b111111111111111111;
        watermark[1262] <= 18'b111000000000000000;
        watermark[1263] <= 18'b000000000000000000;
        watermark[1264] <= 18'b000000000011111111;
        watermark[1265] <= 18'b111111111111111111;
        watermark[1266] <= 18'b111111111111111111;
        watermark[1267] <= 18'b111111111111111111;
        watermark[1268] <= 18'b111111111111111100;
        watermark[1269] <= 18'b000000000000000000;
        watermark[1270] <= 18'b000000000000000000;
        watermark[1271] <= 18'b000011111111111111;
        watermark[1272] <= 18'b111111111111111111;
        watermark[1273] <= 18'b111100000000000000;
        watermark[1274] <= 18'b000000000000000000;
        watermark[1275] <= 18'b000000000011111111;
        watermark[1276] <= 18'b111111111111111111;
        watermark[1277] <= 18'b111111111111111111;
        watermark[1278] <= 18'b111111111111111111;
        watermark[1279] <= 18'b111111111111111111;
        watermark[1280] <= 18'b100000000000000000;
        watermark[1281] <= 18'b000000000000000000;
        watermark[1282] <= 18'b000000001111111111;
        watermark[1283] <= 18'b111111111111111111;
        watermark[1284] <= 18'b111100000000000000;
        watermark[1285] <= 18'b000000000000000000;
        watermark[1286] <= 18'b000000000011111111;
        watermark[1287] <= 18'b111111111111111111;
        watermark[1288] <= 18'b111111111111111111;
        watermark[1289] <= 18'b111111111111111111;
        watermark[1290] <= 18'b111111111111111111;
        watermark[1291] <= 18'b111111000000000000;
        watermark[1292] <= 18'b000000000000000000;
        watermark[1293] <= 18'b000000000001111111;
        watermark[1294] <= 18'b111111111111111111;
        watermark[1295] <= 18'b111110000000000000;
        watermark[1296] <= 18'b000000000000000000;
        watermark[1297] <= 18'b000000000011111111;
        watermark[1298] <= 18'b111111111111111111;
        watermark[1299] <= 18'b111111111111111111;
        watermark[1300] <= 18'b111111111111111111;
        watermark[1301] <= 18'b111111111111111111;
        watermark[1302] <= 18'b111111111110000000;
        watermark[1303] <= 18'b000000000000000000;
        watermark[1304] <= 18'b000000000000001111;
        watermark[1305] <= 18'b111111111111111111;
        watermark[1306] <= 18'b111111000000000000;
        watermark[1307] <= 18'b000000000000000000;
        watermark[1308] <= 18'b000000000111111111;
        watermark[1309] <= 18'b111111111111111111;
        watermark[1310] <= 18'b111111111111111111;
        watermark[1311] <= 18'b111111111111111111;
        watermark[1312] <= 18'b111111111111111111;
        watermark[1313] <= 18'b111111111111111111;
        watermark[1314] <= 18'b111111111111111111;
        watermark[1315] <= 18'b111111111111111111;
        watermark[1316] <= 18'b111111111111111111;
        watermark[1317] <= 18'b111111111111111111;
        watermark[1318] <= 18'b111111111111111111;
        watermark[1319] <= 18'b111111111111111111;
        watermark[1320] <= 18'b111111111111111111;
        watermark[1321] <= 18'b111111111111111111;
        watermark[1322] <= 18'b111111111111111111;
        watermark[1323] <= 18'b111111111111111111;
        watermark[1324] <= 18'b111111111111111111;
        watermark[1325] <= 18'b111111111111111111;
        watermark[1326] <= 18'b111111111111111111;
        watermark[1327] <= 18'b111111111111111111;
        watermark[1328] <= 18'b111111111111111111;
        watermark[1329] <= 18'b111111111111111111;
        watermark[1330] <= 18'b111111111111111111;
        watermark[1331] <= 18'b111111111111111111;
        watermark[1332] <= 18'b111111111111111111;
        watermark[1333] <= 18'b111111111111111111;
        watermark[1334] <= 18'b111111111111111111;
        watermark[1335] <= 18'b111111111111111111;
        watermark[1336] <= 18'b111111111111111111;
        watermark[1337] <= 18'b111111111111111111;
        watermark[1338] <= 18'b111111111111111111;
        watermark[1339] <= 18'b111111111111111111;
        watermark[1340] <= 18'b111111111111111111;
        watermark[1341] <= 18'b111111111111111111;
        watermark[1342] <= 18'b111111111111111111;
        watermark[1343] <= 18'b111111111111111111;
        watermark[1344] <= 18'b111111111111111111;
        watermark[1345] <= 18'b111111111111111111;
        watermark[1346] <= 18'b111111111111111111;
        watermark[1347] <= 18'b111111111111111111;
        watermark[1348] <= 18'b111111111111111111;
        watermark[1349] <= 18'b111111111111111111;
        watermark[1350] <= 18'b111111111111111111;
        watermark[1351] <= 18'b111111111111111111;
        watermark[1352] <= 18'b111111111111111111;
        watermark[1353] <= 18'b111111111111111111;
        watermark[1354] <= 18'b111111111111111111;
        watermark[1355] <= 18'b111111111111111111;
        watermark[1356] <= 18'b111111111111111111;
        watermark[1357] <= 18'b111111111111111111;
        watermark[1358] <= 18'b111111111111000000;
        watermark[1359] <= 18'b000000000000000000;
        watermark[1360] <= 18'b000001111111111111;
        watermark[1361] <= 18'b111111111111111100;
        watermark[1362] <= 18'b000000000000000000;
        watermark[1363] <= 18'b000000000111111111;
        watermark[1364] <= 18'b111111111111111111;
        watermark[1365] <= 18'b111111111111111111;
        watermark[1366] <= 18'b111111111111111111;
        watermark[1367] <= 18'b111111111111111111;
        watermark[1368] <= 18'b111111111111111100;
        watermark[1369] <= 18'b000000000000000000;
        watermark[1370] <= 18'b000000000000000000;
        watermark[1371] <= 18'b000000111111111111;
        watermark[1372] <= 18'b111111111111111111;
        watermark[1373] <= 18'b110000000000000000;
        watermark[1374] <= 18'b000000000000000000;
        watermark[1375] <= 18'b000000000111111111;
        watermark[1376] <= 18'b111111111111111111;
        watermark[1377] <= 18'b111111111111111111;
        watermark[1378] <= 18'b111111111111111111;
        watermark[1379] <= 18'b111111111111111111;
        watermark[1380] <= 18'b100000000000000000;
        watermark[1381] <= 18'b000000000000000000;
        watermark[1382] <= 18'b000000011111111111;
        watermark[1383] <= 18'b111111111111111111;
        watermark[1384] <= 18'b111110000000000000;
        watermark[1385] <= 18'b000000000000000000;
        watermark[1386] <= 18'b000000000001111111;
        watermark[1387] <= 18'b111111111111111111;
        watermark[1388] <= 18'b111111111111111111;
        watermark[1389] <= 18'b111111111111111111;
        watermark[1390] <= 18'b111111111111111111;
        watermark[1391] <= 18'b111100000000000000;
        watermark[1392] <= 18'b000000000000000000;
        watermark[1393] <= 18'b000000011111111111;
        watermark[1394] <= 18'b111111111111111111;
        watermark[1395] <= 18'b111111111000000000;
        watermark[1396] <= 18'b000000000000000000;
        watermark[1397] <= 18'b000000000000111111;
        watermark[1398] <= 18'b111111111111111111;
        watermark[1399] <= 18'b111111111111111111;
        watermark[1400] <= 18'b111111111111111111;
        watermark[1401] <= 18'b111111111111111111;
        watermark[1402] <= 18'b111111000000000000;
        watermark[1403] <= 18'b000000000000000000;
        watermark[1404] <= 18'b000000001111111111;
        watermark[1405] <= 18'b111111111111111111;
        watermark[1406] <= 18'b111111111111000000;
        watermark[1407] <= 18'b000000000000000000;
        watermark[1408] <= 18'b000000000000001111;
        watermark[1409] <= 18'b111111111111111111;
        watermark[1410] <= 18'b111111111111111111;
        watermark[1411] <= 18'b111111111111111111;
        watermark[1412] <= 18'b111111111111111111;
        watermark[1413] <= 18'b111111111000000000;
        watermark[1414] <= 18'b000000000000000000;
        watermark[1415] <= 18'b000000001111111111;
        watermark[1416] <= 18'b111111111111111111;
        watermark[1417] <= 18'b111111111111111000;
        watermark[1418] <= 18'b000000000000000000;
        watermark[1419] <= 18'b000000000000000111;
        watermark[1420] <= 18'b111111111111111111;
        watermark[1421] <= 18'b111111111111111111;
        watermark[1422] <= 18'b111111111111111111;
        watermark[1423] <= 18'b111111111111111111;
        watermark[1424] <= 18'b111111111111000000;
        watermark[1425] <= 18'b000000000000000000;
        watermark[1426] <= 18'b000000000111111111;
        watermark[1427] <= 18'b111111111111111111;
        watermark[1428] <= 18'b111111111111111111;
        watermark[1429] <= 18'b100000000000000000;
        watermark[1430] <= 18'b000000000000000011;
        watermark[1431] <= 18'b111111111111111111;
        watermark[1432] <= 18'b111111111111111111;
        watermark[1433] <= 18'b111111111111111111;
        watermark[1434] <= 18'b111111111111111111;
        watermark[1435] <= 18'b111111111111111000;
        watermark[1436] <= 18'b000000000000000000;
        watermark[1437] <= 18'b000000000111111111;
        watermark[1438] <= 18'b111111111111111111;
        watermark[1439] <= 18'b111111111111111111;
        watermark[1440] <= 18'b111110000000000000;
        watermark[1441] <= 18'b000000000000000001;
        watermark[1442] <= 18'b111111111111111111;
        watermark[1443] <= 18'b111111111111111111;
        watermark[1444] <= 18'b111111111111111111;
        watermark[1445] <= 18'b111111111111111111;
        watermark[1446] <= 18'b111111111111111111;
        watermark[1447] <= 18'b000000000000000000;
        watermark[1448] <= 18'b000000000011111111;
        watermark[1449] <= 18'b111111111111111111;
        watermark[1450] <= 18'b111111111111111111;
        watermark[1451] <= 18'b111111110000000000;
        watermark[1452] <= 18'b000000000000000000;
        watermark[1453] <= 18'b111111111111111111;
        watermark[1454] <= 18'b111111111111111111;
        watermark[1455] <= 18'b111111111111111111;
        watermark[1456] <= 18'b111111111111111111;
        watermark[1457] <= 18'b111111111111111111;
        watermark[1458] <= 18'b111000000000000000;
        watermark[1459] <= 18'b000000000011111111;
        watermark[1460] <= 18'b111111111111111111;
        watermark[1461] <= 18'b111111111111111111;
        watermark[1462] <= 18'b111111111111000000;
        watermark[1463] <= 18'b000000000000000000;
        watermark[1464] <= 18'b011111111111111111;
        watermark[1465] <= 18'b111111111111111111;
        watermark[1466] <= 18'b111111111111111111;
        watermark[1467] <= 18'b111111111111111111;
        watermark[1468] <= 18'b111111111111111111;
        watermark[1469] <= 18'b111111000000000000;
        watermark[1470] <= 18'b000000000011111111;
        watermark[1471] <= 18'b111111111111111111;
        watermark[1472] <= 18'b111111111111111111;
        watermark[1473] <= 18'b111111111111111000;
        watermark[1474] <= 18'b000000000000000000;
        watermark[1475] <= 18'b001111111111111111;
        watermark[1476] <= 18'b111111111111111111;
        watermark[1477] <= 18'b111111111111111111;
        watermark[1478] <= 18'b111111111111111111;
        watermark[1479] <= 18'b111111111111111111;
        watermark[1480] <= 18'b111111111000000000;
        watermark[1481] <= 18'b000000000001111111;
        watermark[1482] <= 18'b111111111111111111;
        watermark[1483] <= 18'b111111111111111111;
        watermark[1484] <= 18'b111111111111111111;
        watermark[1485] <= 18'b100000000000000000;
        watermark[1486] <= 18'b000111111111111111;
        watermark[1487] <= 18'b111111111111111111;
        watermark[1488] <= 18'b111111111111111111;
        watermark[1489] <= 18'b111111111111111111;
        watermark[1490] <= 18'b111111111111111111;
        watermark[1491] <= 18'b111111111111100000;
        watermark[1492] <= 18'b000000000001111111;
        watermark[1493] <= 18'b111111111111111111;
        watermark[1494] <= 18'b111111111111111111;
        watermark[1495] <= 18'b111111111111111111;
        watermark[1496] <= 18'b111110000000000000;
        watermark[1497] <= 18'b000111111111111111;
        watermark[1498] <= 18'b111111111111111111;
        watermark[1499] <= 18'b111111111111111111;
        watermark[1500] <= 18'b111111111111111111;
        watermark[1501] <= 18'b111111111111111111;
        watermark[1502] <= 18'b111111111111111110;
        watermark[1503] <= 18'b000000000001111111;
        watermark[1504] <= 18'b111111111111111111;
        watermark[1505] <= 18'b111111111111111111;
        watermark[1506] <= 18'b111111111111111111;
        watermark[1507] <= 18'b111111111000000000;
        watermark[1508] <= 18'b000111111111111111;
        watermark[1509] <= 18'b111111111111111111;
        watermark[1510] <= 18'b111111111111111111;
        watermark[1511] <= 18'b111111111111111111;
        watermark[1512] <= 18'b111111111111111111;
        watermark[1513] <= 18'b111111111111111111;
        watermark[1514] <= 18'b111000000011111111;
        watermark[1515] <= 18'b111111111111111111;
        watermark[1516] <= 18'b111111111111111111;
        watermark[1517] <= 18'b111111111111111111;
        watermark[1518] <= 18'b111111111111110000;
        watermark[1519] <= 18'b000111111111111111;
        watermark[1520] <= 18'b111111111111111111;
        watermark[1521] <= 18'b111111111111111111;
        watermark[1522] <= 18'b111111111111111111;
        watermark[1523] <= 18'b111111111111111111;
        watermark[1524] <= 18'b111111111111111111;
        watermark[1525] <= 18'b111111111111111111;
        watermark[1526] <= 18'b111111111111111111;
        watermark[1527] <= 18'b111111111111111111;
        watermark[1528] <= 18'b111111111111111111;
        watermark[1529] <= 18'b111111111111111111;
        watermark[1530] <= 18'b111111111111111111;
        watermark[1531] <= 18'b111111111111111111;
        watermark[1532] <= 18'b111111111111111111;
        watermark[1533] <= 18'b111111111111111111;
        watermark[1534] <= 18'b111111111111111111;
        watermark[1535] <= 18'b111111111111111111;
        watermark[1536] <= 18'b111111111111111111;
        watermark[1537] <= 18'b111111111111111111;
        watermark[1538] <= 18'b111111111111111111;
        watermark[1539] <= 18'b111111111111111111;
        watermark[1540] <= 18'b111111111111111111;
        watermark[1541] <= 18'b111111111111111111;
        watermark[1542] <= 18'b111111111111111111;
        watermark[1543] <= 18'b111111111111111111;
        watermark[1544] <= 18'b111111111111111111;
        watermark[1545] <= 18'b111111111111111111;
        watermark[1546] <= 18'b111111111111111111;
        watermark[1547] <= 18'b111111111111111111;
        watermark[1548] <= 18'b111111111111111111;
        watermark[1549] <= 18'b111111111111111111;
        watermark[1550] <= 18'b111111111111111111;
        watermark[1551] <= 18'b111111111111111111;
        watermark[1552] <= 18'b111111111111111111;
        watermark[1553] <= 18'b111111111111111111;
        watermark[1554] <= 18'b111111111111111111;
        watermark[1555] <= 18'b111111111111111111;
        watermark[1556] <= 18'b111111111111111111;
        watermark[1557] <= 18'b111111111111111111;
        watermark[1558] <= 18'b111111111111111111;
        watermark[1559] <= 18'b111111111111111111;
        watermark[1560] <= 18'b111111111111111111;
        watermark[1561] <= 18'b111111111111111111;
        watermark[1562] <= 18'b111111111111111111;
        watermark[1563] <= 18'b111111111111111111;
        watermark[1564] <= 18'b111111111111111111;
        watermark[1565] <= 18'b111111111111111111;
        watermark[1566] <= 18'b111111111111111111;
        watermark[1567] <= 18'b111111111111111111;
        watermark[1568] <= 18'b111111111111111111;
        watermark[1569] <= 18'b111111111111111111;
        watermark[1570] <= 18'b111111111111111111;
        watermark[1571] <= 18'b111111111111111111;
        watermark[1572] <= 18'b111111111111111111;
        watermark[1573] <= 18'b111111111111111111;
        watermark[1574] <= 18'b111111111111111111;
        watermark[1575] <= 18'b111111111111111111;
        watermark[1576] <= 18'b111111111111111111;
        watermark[1577] <= 18'b111111111111111111;
        watermark[1578] <= 18'b111111111111111111;
        watermark[1579] <= 18'b111111111111111111;
        watermark[1580] <= 18'b111111111111111111;
        watermark[1581] <= 18'b111111111111111111;
        watermark[1582] <= 18'b111111111111111111;
        watermark[1583] <= 18'b111111111111111111;
        watermark[1584] <= 18'b111111111111111111;
        watermark[1585] <= 18'b111111111111111111;
        watermark[1586] <= 18'b111111111111111111;
        watermark[1587] <= 18'b111111111111111111;
        watermark[1588] <= 18'b111111111111111111;
        watermark[1589] <= 18'b111111111111111111;
        watermark[1590] <= 18'b111111111111111111;
        watermark[1591] <= 18'b111111111111111111;
        watermark[1592] <= 18'b111111111111111111;
        watermark[1593] <= 18'b111111111111111111;
        watermark[1594] <= 18'b111111111111111111;
        watermark[1595] <= 18'b111111111111111111;
        watermark[1596] <= 18'b111111111111111111;
        watermark[1597] <= 18'b111111111111111111;
        watermark[1598] <= 18'b111111111111111111;
        watermark[1599] <= 18'b111111111111111111;
        watermark[1600] <= 18'b111111111111111111;
        watermark[1601] <= 18'b111111111111111111;
        watermark[1602] <= 18'b111111111111111111;
        watermark[1603] <= 18'b111111111111111111;
        watermark[1604] <= 18'b111111111111111111;
        watermark[1605] <= 18'b111111111111111111;
        watermark[1606] <= 18'b111111111111111111;
        watermark[1607] <= 18'b111111111111111111;
        watermark[1608] <= 18'b111111111111111111;
        watermark[1609] <= 18'b111111111111111111;
        watermark[1610] <= 18'b111111111111111111;
        watermark[1611] <= 18'b111111111111111111;
        watermark[1612] <= 18'b111111111111111111;
        watermark[1613] <= 18'b111111111111111111;
        watermark[1614] <= 18'b111111111111111111;
        watermark[1615] <= 18'b111111111111111111;
        watermark[1616] <= 18'b111111111111111111;
        watermark[1617] <= 18'b111111111111111111;
        watermark[1618] <= 18'b111111111111111111;
        watermark[1619] <= 18'b111111111111111111;
        watermark[1620] <= 18'b111111111111111111;
        watermark[1621] <= 18'b111111111111111111;
        watermark[1622] <= 18'b111111111111111111;
        watermark[1623] <= 18'b111111111111111111;
        watermark[1624] <= 18'b111111111111111111;
        watermark[1625] <= 18'b111111111111111111;
        watermark[1626] <= 18'b111111111111111111;
        watermark[1627] <= 18'b111111111111111111;
        watermark[1628] <= 18'b111111111111111111;
        watermark[1629] <= 18'b111111111111111111;
        watermark[1630] <= 18'b111111111111111111;
        watermark[1631] <= 18'b111111111111111111;
        watermark[1632] <= 18'b111111111111111111;
        watermark[1633] <= 18'b111111111111111111;
        watermark[1634] <= 18'b111111111111111111;
        watermark[1635] <= 18'b111111111111111111;
        watermark[1636] <= 18'b111111111111111111;
        watermark[1637] <= 18'b111111111111111111;
        watermark[1638] <= 18'b111111111111111111;
        watermark[1639] <= 18'b111111111111111111;
        watermark[1640] <= 18'b111111111111111111;
        watermark[1641] <= 18'b111111111111111111;
        watermark[1642] <= 18'b111111111111111111;
        watermark[1643] <= 18'b111111111111111111;
        watermark[1644] <= 18'b111111111111111111;
        watermark[1645] <= 18'b111111111111111111;
        watermark[1646] <= 18'b111111111111111111;
        watermark[1647] <= 18'b111111111111111111;
        watermark[1648] <= 18'b111111111111111111;
        watermark[1649] <= 18'b111111111111111111;
        watermark[1650] <= 18'b111111111111111111;
        watermark[1651] <= 18'b111111111111111111;
        watermark[1652] <= 18'b111111111111111111;
        watermark[1653] <= 18'b111111111111111111;
        watermark[1654] <= 18'b111111111111111111;
        watermark[1655] <= 18'b111111111111111111;
        watermark[1656] <= 18'b111111111111111111;
        watermark[1657] <= 18'b100000111111111111;
        watermark[1658] <= 18'b000000111100000111;
        watermark[1659] <= 18'b111111111000001111;
        watermark[1660] <= 18'b111111110000001111;
        watermark[1661] <= 18'b111000000111111111;
        watermark[1662] <= 18'b110000001111111111;
        watermark[1663] <= 18'b100000111111111100;
        watermark[1664] <= 18'b000000000001111000;
        watermark[1665] <= 18'b000111111111111111;
        watermark[1666] <= 18'b111111111111111111;
        watermark[1667] <= 18'b111111111111111111;
        watermark[1668] <= 18'b111000001111111111;
        watermark[1669] <= 18'b110000001111000001;
        watermark[1670] <= 18'b111111111110000011;
        watermark[1671] <= 18'b111111111000000011;
        watermark[1672] <= 18'b111111000001111111;
        watermark[1673] <= 18'b111000000011111111;
        watermark[1674] <= 18'b111000001111111000;
        watermark[1675] <= 18'b000000000000011110;
        watermark[1676] <= 18'b000001111111111111;
        watermark[1677] <= 18'b111111111111111111;
        watermark[1678] <= 18'b111111111111111111;
        watermark[1679] <= 18'b111110000011111111;
        watermark[1680] <= 18'b111100000011110000;
        watermark[1681] <= 18'b011111111111100000;
        watermark[1682] <= 18'b111111111110000000;
        watermark[1683] <= 18'b011111110000001111;
        watermark[1684] <= 18'b111110000000011111;
        watermark[1685] <= 18'b111100000011111100;
        watermark[1686] <= 18'b000000000000000111;
        watermark[1687] <= 18'b100000011111111111;
        watermark[1688] <= 18'b111111111111111111;
        watermark[1689] <= 18'b111111111111111111;
        watermark[1690] <= 18'b111111100000111111;
        watermark[1691] <= 18'b111111000000111100;
        watermark[1692] <= 18'b000111111111111000;
        watermark[1693] <= 18'b001111111111000000;
        watermark[1694] <= 18'b000111111100000011;
        watermark[1695] <= 18'b111111100000000111;
        watermark[1696] <= 18'b111111000000111100;
        watermark[1697] <= 18'b000000000000000001;
        watermark[1698] <= 18'b111000000111111111;
        watermark[1699] <= 18'b111111111111111111;
        watermark[1700] <= 18'b111111111111111111;
        watermark[1701] <= 18'b111111111000001111;
        watermark[1702] <= 18'b111111110000001111;
        watermark[1703] <= 18'b000001111111111110;
        watermark[1704] <= 18'b000011111111110000;
        watermark[1705] <= 18'b000000111111100000;
        watermark[1706] <= 18'b111111110000000001;
        watermark[1707] <= 18'b111111110000011111;
        watermark[1708] <= 18'b000000000111111111;
        watermark[1709] <= 18'b111110000001111111;
        watermark[1710] <= 18'b111111111111111111;
        watermark[1711] <= 18'b111111111111111111;
        watermark[1712] <= 18'b111111111110000011;
        watermark[1713] <= 18'b111111111100000011;
        watermark[1714] <= 18'b110000011111111111;
        watermark[1715] <= 18'b100000111111111000;
        watermark[1716] <= 18'b000000001111111000;
        watermark[1717] <= 18'b000111111100000000;
        watermark[1718] <= 18'b001111111100000111;
        watermark[1719] <= 18'b100000001111111111;
        watermark[1720] <= 18'b111111100000011111;
        watermark[1721] <= 18'b111111111111111111;
        watermark[1722] <= 18'b111111111111111111;
        watermark[1723] <= 18'b111111111111100000;
        watermark[1724] <= 18'b111111111111000000;
        watermark[1725] <= 18'b111100000111111111;
        watermark[1726] <= 18'b111000001111111110;
        watermark[1727] <= 18'b000010000001111110;
        watermark[1728] <= 18'b000001111111000000;
        watermark[1729] <= 18'b000011111110000001;
        watermark[1730] <= 18'b111000000111111111;
        watermark[1731] <= 18'b111111111000000111;
        watermark[1732] <= 18'b111111111111111111;
        watermark[1733] <= 18'b111111111111111111;
        watermark[1734] <= 18'b111111111111111000;
        watermark[1735] <= 18'b001111111111110000;
        watermark[1736] <= 18'b001111000001111111;
        watermark[1737] <= 18'b111110000011111111;
        watermark[1738] <= 18'b100000110000011111;
        watermark[1739] <= 18'b110000011111110000;
        watermark[1740] <= 18'b000000111111100000;
        watermark[1741] <= 18'b111100000011111111;
        watermark[1742] <= 18'b111111111110000001;
        watermark[1743] <= 18'b111111111111111111;
        watermark[1744] <= 18'b111111111111111111;
        watermark[1745] <= 18'b111111111111111110;
        watermark[1746] <= 18'b000011111111111100;
        watermark[1747] <= 18'b000011110000011111;
        watermark[1748] <= 18'b111111100000111111;
        watermark[1749] <= 18'b110000011100000111;
        watermark[1750] <= 18'b111100000011111000;
        watermark[1751] <= 18'b001000000111111000;
        watermark[1752] <= 18'b001111000000111111;
        watermark[1753] <= 18'b111111111111100000;
        watermark[1754] <= 18'b011111111111111111;
        watermark[1755] <= 18'b111111111111111111;
        watermark[1756] <= 18'b111111111111111111;
        watermark[1757] <= 18'b100000011111111111;
        watermark[1758] <= 18'b000000111100000111;
        watermark[1759] <= 18'b111111111000001111;
        watermark[1760] <= 18'b111100000111000000;
        watermark[1761] <= 18'b111111000000111110;
        watermark[1762] <= 18'b000011000001111100;
        watermark[1763] <= 18'b000011110000001111;
        watermark[1764] <= 18'b111111111111111000;
        watermark[1765] <= 18'b000111111111111111;
        watermark[1766] <= 18'b111111111111111111;
        watermark[1767] <= 18'b111111111111111111;
        watermark[1768] <= 18'b111000000000000000;
        watermark[1769] <= 18'b000000001111000001;
        watermark[1770] <= 18'b111111111110000011;
        watermark[1771] <= 18'b111110000011111000;
        watermark[1772] <= 18'b001111111000001111;
        watermark[1773] <= 18'b100000110000011111;
        watermark[1774] <= 18'b000001111100000000;
        watermark[1775] <= 18'b000000000000011110;
        watermark[1776] <= 18'b000001111111111111;
        watermark[1777] <= 18'b111111111111111111;
        watermark[1778] <= 18'b111111111111111111;
        watermark[1779] <= 18'b111110000000000000;
        watermark[1780] <= 18'b000000000011110000;
        watermark[1781] <= 18'b011111111111100000;
        watermark[1782] <= 18'b111111100000111110;
        watermark[1783] <= 18'b000001111110000001;
        watermark[1784] <= 18'b111000001100000011;
        watermark[1785] <= 18'b110000011111000000;
        watermark[1786] <= 18'b000000000000000111;
        watermark[1787] <= 18'b100000011111111111;
        watermark[1788] <= 18'b111111111111111111;
        watermark[1789] <= 18'b111111111111111111;
        watermark[1790] <= 18'b111111100000000000;
        watermark[1791] <= 18'b000000000000111100;
        watermark[1792] <= 18'b000111111111111000;
        watermark[1793] <= 18'b001111110000001111;
        watermark[1794] <= 18'b110000011111100000;
        watermark[1795] <= 18'b011100000111100000;
        watermark[1796] <= 18'b111000000111110000;
        watermark[1797] <= 18'b000000000000000001;
        watermark[1798] <= 18'b111000000111111111;
        watermark[1799] <= 18'b111111111111111111;
        watermark[1800] <= 18'b111111111111111111;
        watermark[1801] <= 18'b111111111000000000;
        watermark[1802] <= 18'b000000000000001111;
        watermark[1803] <= 18'b000001111111111110;
        watermark[1804] <= 18'b000011111100000111;
        watermark[1805] <= 18'b111100000011111100;
        watermark[1806] <= 18'b000111000001111000;
        watermark[1807] <= 18'b001110000011111100;
        watermark[1808] <= 18'b000000000000000000;
        watermark[1809] <= 18'b011110000001111111;
        watermark[1810] <= 18'b111111111111111111;
        watermark[1811] <= 18'b111111111111111111;
        watermark[1812] <= 18'b111111111110000011;
        watermark[1813] <= 18'b111111111100000011;
        watermark[1814] <= 18'b110000011111111111;
        watermark[1815] <= 18'b100000111110000000;
        watermark[1816] <= 18'b000000000000111111;
        watermark[1817] <= 18'b000000110000011110;
        watermark[1818] <= 18'b000001100000111111;
        watermark[1819] <= 18'b000000111111111111;
        watermark[1820] <= 18'b111111100000011111;
        watermark[1821] <= 18'b111111111111111111;
        watermark[1822] <= 18'b111111111111111111;
        watermark[1823] <= 18'b111111111111100000;
        watermark[1824] <= 18'b111111111111000000;
        watermark[1825] <= 18'b111100000111111111;
        watermark[1826] <= 18'b111000001111100000;
        watermark[1827] <= 18'b000000000000000111;
        watermark[1828] <= 18'b111000001000001111;
        watermark[1829] <= 18'b110000011000001111;
        watermark[1830] <= 18'b110000001111111111;
        watermark[1831] <= 18'b111111111000000111;
        watermark[1832] <= 18'b111111111111111111;
        watermark[1833] <= 18'b111111111111111111;
        watermark[1834] <= 18'b111111111111111000;
        watermark[1835] <= 18'b001111111111110000;
        watermark[1836] <= 18'b001111000000111111;
        watermark[1837] <= 18'b111110000011110000;
        watermark[1838] <= 18'b000000000000000001;
        watermark[1839] <= 18'b111110000010000011;
        watermark[1840] <= 18'b111100000100000111;
        watermark[1841] <= 18'b111100000011111111;
        watermark[1842] <= 18'b111111111110000001;
        watermark[1843] <= 18'b111111111111111111;
        watermark[1844] <= 18'b111111111111111111;
        watermark[1845] <= 18'b111111111111111110;
        watermark[1846] <= 18'b000011111111111100;
        watermark[1847] <= 18'b000011110000001111;
        watermark[1848] <= 18'b111111000000111100;
        watermark[1849] <= 18'b000000000000000000;
        watermark[1850] <= 18'b001111100000000000;
        watermark[1851] <= 18'b111111000000000001;
        watermark[1852] <= 18'b111111100000011111;
        watermark[1853] <= 18'b111111111111100000;
        watermark[1854] <= 18'b011111111111111111;
        watermark[1855] <= 18'b111111111111111111;
        watermark[1856] <= 18'b111111111111111111;
        watermark[1857] <= 18'b100000111111111111;
        watermark[1858] <= 18'b000000111100000011;
        watermark[1859] <= 18'b111111110000001111;
        watermark[1860] <= 18'b000001111111111100;
        watermark[1861] <= 18'b000011111100000000;
        watermark[1862] <= 18'b001111111000000000;
        watermark[1863] <= 18'b011111111000000011;
        watermark[1864] <= 18'b111111111111111000;
        watermark[1865] <= 18'b000111111111111111;
        watermark[1866] <= 18'b111111111111111111;
        watermark[1867] <= 18'b111111111111111111;
        watermark[1868] <= 18'b111000001111111111;
        watermark[1869] <= 18'b110000001111100000;
        watermark[1870] <= 18'b001111111000000111;
        watermark[1871] <= 18'b100000011111111111;
        watermark[1872] <= 18'b100000011111000000;
        watermark[1873] <= 18'b000111111110000000;
        watermark[1874] <= 18'b001111111111000000;
        watermark[1875] <= 18'b001111111111111110;
        watermark[1876] <= 18'b000001111111111111;
        watermark[1877] <= 18'b111111111111111111;
        watermark[1878] <= 18'b111111111111111111;
        watermark[1879] <= 18'b111110000011111111;
        watermark[1880] <= 18'b111100000011111000;
        watermark[1881] <= 18'b000000000000000001;
        watermark[1882] <= 18'b111000001111111111;
        watermark[1883] <= 18'b111000000111110000;
        watermark[1884] <= 18'b000001111111100000;
        watermark[1885] <= 18'b000011111111110000;
        watermark[1886] <= 18'b000000000000000111;
        watermark[1887] <= 18'b100000011111111111;
        watermark[1888] <= 18'b111111111111111111;
        watermark[1889] <= 18'b111111111111111111;
        watermark[1890] <= 18'b111111100000111111;
        watermark[1891] <= 18'b111111000000111111;
        watermark[1892] <= 18'b000000000000000000;
        watermark[1893] <= 18'b111100000011111111;
        watermark[1894] <= 18'b111110000001111110;
        watermark[1895] <= 18'b000000011111111100;
        watermark[1896] <= 18'b000000111111111110;
        watermark[1897] <= 18'b000000000000000001;
        watermark[1898] <= 18'b111000000111111111;
        watermark[1899] <= 18'b111111111111111111;
        watermark[1900] <= 18'b111111111111111111;
        watermark[1901] <= 18'b111111111000001111;
        watermark[1902] <= 18'b111111110000001111;
        watermark[1903] <= 18'b111100000000000000;
        watermark[1904] <= 18'b011111000001111111;
        watermark[1905] <= 18'b111111110000001111;
        watermark[1906] <= 18'b100000000111111111;
        watermark[1907] <= 18'b000000011111111111;
        watermark[1908] <= 18'b111000000000000000;
        watermark[1909] <= 18'b011110000001111111;
        watermark[1910] <= 18'b111111111111111111;
        watermark[1911] <= 18'b111111111111111111;
        watermark[1912] <= 18'b111111111110000011;
        watermark[1913] <= 18'b111111111100000011;
        watermark[1914] <= 18'b111111110000000000;
        watermark[1915] <= 18'b111111100000011111;
        watermark[1916] <= 18'b111111111100000011;
        watermark[1917] <= 18'b111100000011111111;
        watermark[1918] <= 18'b110000000111111111;
        watermark[1919] <= 18'b111111110000000000;
        watermark[1920] <= 18'b000111100000011111;
        watermark[1921] <= 18'b111111111111111111;
        watermark[1922] <= 18'b111111111111111111;
        watermark[1923] <= 18'b111111111111111111;
        watermark[1924] <= 18'b111111111111111111;
        watermark[1925] <= 18'b111111111111111111;
        watermark[1926] <= 18'b111111111111111111;
        watermark[1927] <= 18'b111111111111111111;
        watermark[1928] <= 18'b111111111111111111;
        watermark[1929] <= 18'b111111111111111111;
        watermark[1930] <= 18'b111111111111111111;
        watermark[1931] <= 18'b111111111111111111;
        watermark[1932] <= 18'b111111111111111111;
        watermark[1933] <= 18'b111111111111111111;
        watermark[1934] <= 18'b111111111111111111;
        watermark[1935] <= 18'b111111111111111111;
        watermark[1936] <= 18'b111111111111111111;
        watermark[1937] <= 18'b111111111111111111;
        watermark[1938] <= 18'b111111111111111111;
        watermark[1939] <= 18'b111111111111111111;
        watermark[1940] <= 18'b111111111111111111;
        watermark[1941] <= 18'b111111111111111111;
        watermark[1942] <= 18'b111111111111111111;
        watermark[1943] <= 18'b111111111111111111;
        watermark[1944] <= 18'b111111111111111111;
        watermark[1945] <= 18'b111111111111111111;
        watermark[1946] <= 18'b111111111111111111;
        watermark[1947] <= 18'b111111111111111111;
        watermark[1948] <= 18'b111111111111111111;
        watermark[1949] <= 18'b111111111111111111;
        watermark[1950] <= 18'b111111111111111111;
        watermark[1951] <= 18'b111111111111111111;
        watermark[1952] <= 18'b111111111111111111;
        watermark[1953] <= 18'b111111111111111111;
        watermark[1954] <= 18'b111111111111111111;
        watermark[1955] <= 18'b111111111111111111;
        watermark[1956] <= 18'b111111111111111111;
        watermark[1957] <= 18'b111111111111111111;
        watermark[1958] <= 18'b111111111111111111;
        watermark[1959] <= 18'b111111111111111111;
        watermark[1960] <= 18'b111111111111111111;
        watermark[1961] <= 18'b111111111111111111;
        watermark[1962] <= 18'b111111111111111111;
        watermark[1963] <= 18'b111111111111111111;
        watermark[1964] <= 18'b111111111111111111;
        watermark[1965] <= 18'b111111111111111111;
        watermark[1966] <= 18'b111111111111111111;
        watermark[1967] <= 18'b111111111111111111;
        watermark[1968] <= 18'b111111111111111111;
        watermark[1969] <= 18'b111111111111111111;
        watermark[1970] <= 18'b111111111111111111;
        watermark[1971] <= 18'b111111111111111111;
        watermark[1972] <= 18'b111111111111111111;
        watermark[1973] <= 18'b111111111111111111;
        watermark[1974] <= 18'b111111111111111111;
        watermark[1975] <= 18'b111111111111111111;
        watermark[1976] <= 18'b111111111111111111;
        watermark[1977] <= 18'b111111111111111111;
        watermark[1978] <= 18'b111111111111111111;
        watermark[1979] <= 18'b111111111111111111;
        watermark[1980] <= 18'b111111111111111111;
        watermark[1981] <= 18'b111111111111111111;
        watermark[1982] <= 18'b111111111111111111;
        watermark[1983] <= 18'b111111111111111111;
        watermark[1984] <= 18'b111111111111111111;
        watermark[1985] <= 18'b111111111111111111;
        watermark[1986] <= 18'b111111111111111111;
        watermark[1987] <= 18'b111111111111111111;
        watermark[1988] <= 18'b111111111111111111;
        watermark[1989] <= 18'b111111111111111111;
        watermark[1990] <= 18'b111111111111111111;
        watermark[1991] <= 18'b111111111111111111;
        watermark[1992] <= 18'b111111111111111111;
        watermark[1993] <= 18'b111111111111111111;
        watermark[1994] <= 18'b111111111111111111;
        watermark[1995] <= 18'b111111111111111111;
        watermark[1996] <= 18'b111111111111111111;
        watermark[1997] <= 18'b111111111111111111;
        watermark[1998] <= 18'b111111111111111111;
        watermark[1999] <= 18'b111111111111111111;
        watermark[2000] <= 18'b111111111111111111;
        watermark[2001] <= 18'b111111111111111111;
        watermark[2002] <= 18'b111111111111111111;
        watermark[2003] <= 18'b111111111111111111;
        watermark[2004] <= 18'b111111111111111111;
        watermark[2005] <= 18'b111111111111111111;
        watermark[2006] <= 18'b111111111111111111;
        watermark[2007] <= 18'b111111111111111111;
        watermark[2008] <= 18'b111111111111111111;
        watermark[2009] <= 18'b111111111111111111;
        watermark[2010] <= 18'b111111111111111111;
        watermark[2011] <= 18'b111111111111111111;
        watermark[2012] <= 18'b111111111111111111;
        watermark[2013] <= 18'b111111111111111111;
        watermark[2014] <= 18'b111111111111111111;
        watermark[2015] <= 18'b111111111111111111;
        watermark[2016] <= 18'b111111111111111111;
        watermark[2017] <= 18'b111111111111111111;
        watermark[2018] <= 18'b111111111111111111;
        watermark[2019] <= 18'b111111111111111111;
        watermark[2020] <= 18'b111111111111111111;
        watermark[2021] <= 18'b111111111111111111;
        watermark[2022] <= 18'b111111111111111111;
        watermark[2023] <= 18'b111111111111111111;
        watermark[2024] <= 18'b111111111111111111;
        watermark[2025] <= 18'b111111111111111111;
        watermark[2026] <= 18'b111111111111111111;
        watermark[2027] <= 18'b111111111111111111;
        watermark[2028] <= 18'b111111111111111111;
        watermark[2029] <= 18'b111111111111111111;
        watermark[2030] <= 18'b111111111111111111;
        watermark[2031] <= 18'b111111111111111111;
        watermark[2032] <= 18'b111111111111111111;
        watermark[2033] <= 18'b111111111111111111;
        watermark[2034] <= 18'b111111111111111111;
        watermark[2035] <= 18'b111111111111111111;
        watermark[2036] <= 18'b111111111111111111;
        watermark[2037] <= 18'b111111111111111111;
        watermark[2038] <= 18'b111111111111111111;
        watermark[2039] <= 18'b111111111111111111;
        watermark[2040] <= 18'b111111111111111111;
        watermark[2041] <= 18'b111111111111111111;
        watermark[2042] <= 18'b111111111111111111;
        watermark[2043] <= 18'b111111111111111111;
        watermark[2044] <= 18'b111111111111111111;
        watermark[2045] <= 18'b111111111111111111;
        watermark[2046] <= 18'b111111111111111111;
        watermark[2047] <= 18'b111111111111111111;
        watermark[2048] <= 18'b111111111111111111;
        watermark[2049] <= 18'b111111111111111111;
        watermark[2050] <= 18'b111111111111111111;
        watermark[2051] <= 18'b111111111111111111;
        watermark[2052] <= 18'b111111111111111111;
        watermark[2053] <= 18'b111111111111111111;
        watermark[2054] <= 18'b111111111111111111;
        watermark[2055] <= 18'b111111111111111111;
        watermark[2056] <= 18'b111111111111111111;
        watermark[2057] <= 18'b111111111111111111;
        watermark[2058] <= 18'b111111111111111111;
        watermark[2059] <= 18'b111111111111111111;
        watermark[2060] <= 18'b111111111111111111;
        watermark[2061] <= 18'b111111111111111111;
        watermark[2062] <= 18'b111111111111111111;
        watermark[2063] <= 18'b111111111111111111;
        watermark[2064] <= 18'b111111111111111111;
        watermark[2065] <= 18'b111111111111111111;
        watermark[2066] <= 18'b111111111111111111;
        watermark[2067] <= 18'b111111111111111111;
        watermark[2068] <= 18'b111111111111111111;
        watermark[2069] <= 18'b111111111111111111;
        watermark[2070] <= 18'b111111111111111111;
        watermark[2071] <= 18'b111111111111111111;
        watermark[2072] <= 18'b111111111111111111;
        watermark[2073] <= 18'b111111111111111111;
        watermark[2074] <= 18'b111111111111111111;
        watermark[2075] <= 18'b111111111111111111;
        watermark[2076] <= 18'b111111111111111111;
        watermark[2077] <= 18'b111111111111111111;
        watermark[2078] <= 18'b111111111111111111;
        watermark[2079] <= 18'b111111111111111111;
        watermark[2080] <= 18'b111111111111111111;
        watermark[2081] <= 18'b111111111111111111;
        watermark[2082] <= 18'b111111111111111111;
        watermark[2083] <= 18'b111111111111111111;
        watermark[2084] <= 18'b111111111111111111;
        watermark[2085] <= 18'b111111111111111111;
        watermark[2086] <= 18'b111111111111111111;
        watermark[2087] <= 18'b111111111111111111;
        watermark[2088] <= 18'b111111111111111111;
        watermark[2089] <= 18'b111111111111111111;
        watermark[2090] <= 18'b111111111111111111;
        watermark[2091] <= 18'b111111111111111111;
        watermark[2092] <= 18'b111111111111111111;
        watermark[2093] <= 18'b111111111111111111;
        watermark[2094] <= 18'b111111111111111111;
        watermark[2095] <= 18'b111111111111111111;
        watermark[2096] <= 18'b111111111111111111;
        watermark[2097] <= 18'b111111111111111111;
        watermark[2098] <= 18'b111111111111111111;
        watermark[2099] <= 18'b111111111111111111;
        watermark[2100] <= 18'b111111111111111111;
        watermark[2101] <= 18'b111111111111111111;
        watermark[2102] <= 18'b111111111111111111;
        watermark[2103] <= 18'b111111111111111111;
        watermark[2104] <= 18'b111111111111111111;
        watermark[2105] <= 18'b111111111111111111;
        watermark[2106] <= 18'b111111111111111111;
        watermark[2107] <= 18'b111111111111111111;
        watermark[2108] <= 18'b111111111111111111;
        watermark[2109] <= 18'b111111111111111111;
        watermark[2110] <= 18'b111111111111111111;
        watermark[2111] <= 18'b111111111111111111;
        watermark[2112] <= 18'b111111111111111111;
        watermark[2113] <= 18'b111111111111111111;
        watermark[2114] <= 18'b111111111111111111;
        watermark[2115] <= 18'b111111111111111111;
        watermark[2116] <= 18'b111111111111111111;
        watermark[2117] <= 18'b111111111111111111;
        watermark[2118] <= 18'b111111111111111111;
        watermark[2119] <= 18'b111111111111111111;
        watermark[2120] <= 18'b111111111111111111;
        watermark[2121] <= 18'b111111111111111111;
        watermark[2122] <= 18'b111111111111111111;
        watermark[2123] <= 18'b111111111111111111;
        watermark[2124] <= 18'b111111111111111111;
        watermark[2125] <= 18'b111111111111111111;
        watermark[2126] <= 18'b111111111111111111;
        watermark[2127] <= 18'b111111111111111111;
        watermark[2128] <= 18'b111111111111111111;
        watermark[2129] <= 18'b111111111111111111;
        watermark[2130] <= 18'b111111111111111111;
        watermark[2131] <= 18'b111111111111111111;
        watermark[2132] <= 18'b111111111111111111;
        watermark[2133] <= 18'b111111111111111111;
        watermark[2134] <= 18'b111111111111111111;
        watermark[2135] <= 18'b111111111111111111;
        watermark[2136] <= 18'b111111111111111111;
        watermark[2137] <= 18'b111111111111111111;
        watermark[2138] <= 18'b111111111111111111;
        watermark[2139] <= 18'b111111111111111111;
        watermark[2140] <= 18'b111111111111111111;
        watermark[2141] <= 18'b111111111111111111;
        watermark[2142] <= 18'b111111111111111111;
        watermark[2143] <= 18'b111111111111111111;
        watermark[2144] <= 18'b111111111111111111;
        watermark[2145] <= 18'b111111111111111111;
        watermark[2146] <= 18'b111111111111111111;
        watermark[2147] <= 18'b111111111111111111;
        watermark[2148] <= 18'b111111111111111111;
        watermark[2149] <= 18'b111111111111111111;
        watermark[2150] <= 18'b111111111111111111;
        watermark[2151] <= 18'b111111111111111111;
        watermark[2152] <= 18'b111111111111111111;
        watermark[2153] <= 18'b111111111111111111;
        watermark[2154] <= 18'b111111111111111111;
        watermark[2155] <= 18'b111111111111111111;
        watermark[2156] <= 18'b111111111111111111;
        watermark[2157] <= 18'b111111111111111111;
        watermark[2158] <= 18'b111111111111111111;
        watermark[2159] <= 18'b111111111111111111;
        watermark[2160] <= 18'b111111111111111111;
        watermark[2161] <= 18'b111111111111111111;
        watermark[2162] <= 18'b111111111111111111;
        watermark[2163] <= 18'b111111111111111111;
        watermark[2164] <= 18'b111111111111111111;
        watermark[2165] <= 18'b111111111111111111;
        watermark[2166] <= 18'b111111111111111111;
        watermark[2167] <= 18'b111111111111111111;
        watermark[2168] <= 18'b111111111111111111;
        watermark[2169] <= 18'b111111111111111111;
        watermark[2170] <= 18'b111111111111111111;
        watermark[2171] <= 18'b111111111111111111;
        watermark[2172] <= 18'b111111111111111111;
        watermark[2173] <= 18'b111111111111111111;
        watermark[2174] <= 18'b111111111111111111;
        watermark[2175] <= 18'b111111111111111111;
        watermark[2176] <= 18'b111111111111111111;
        watermark[2177] <= 18'b111111111111111111;
        watermark[2178] <= 18'b111111111111111111;
        watermark[2179] <= 18'b111111111111111111;
        watermark[2180] <= 18'b111111111111111111;
        watermark[2181] <= 18'b111111111111111111;
        watermark[2182] <= 18'b111111111111111111;
        watermark[2183] <= 18'b111111111111111111;
        watermark[2184] <= 18'b111111111111111111;
        watermark[2185] <= 18'b111111111111111111;
        watermark[2186] <= 18'b111111111111111111;
        watermark[2187] <= 18'b111111111111111111;
        watermark[2188] <= 18'b111111111111111111;
        watermark[2189] <= 18'b111111111111111111;
        watermark[2190] <= 18'b111111111111111111;
        watermark[2191] <= 18'b111111111111111111;
        watermark[2192] <= 18'b111111111111111111;
        watermark[2193] <= 18'b111111111111111111;
        watermark[2194] <= 18'b111111111111111111;
        watermark[2195] <= 18'b111111111111111111;
        watermark[2196] <= 18'b111111111111111111;
        watermark[2197] <= 18'b111111111111111111;
        watermark[2198] <= 18'b111111111111111111;
        watermark[2199] <= 18'b111111111111111111;
        watermark[2200] <= 18'b111111111111111111;
        watermark[2201] <= 18'b111111111111111111;
        watermark[2202] <= 18'b111111111111111111;
        watermark[2203] <= 18'b111111111111111111;
        watermark[2204] <= 18'b111111111111111111;
        watermark[2205] <= 18'b111111111111111111;
        watermark[2206] <= 18'b111111111111111111;
        watermark[2207] <= 18'b111111111111111111;
        watermark[2208] <= 18'b111111111111111111;
        watermark[2209] <= 18'b111111111111111111;
        watermark[2210] <= 18'b111111111111111111;
        watermark[2211] <= 18'b111111111111111111;
        watermark[2212] <= 18'b111111111111111111;
        watermark[2213] <= 18'b111111111111111111;
        watermark[2214] <= 18'b111111111111111111;
        watermark[2215] <= 18'b111111111111111111;
        watermark[2216] <= 18'b111111111111111111;
        watermark[2217] <= 18'b111111111111111111;
        watermark[2218] <= 18'b111111111111111111;
        watermark[2219] <= 18'b111111111111111111;
        watermark[2220] <= 18'b111111111111111111;
        watermark[2221] <= 18'b111111111111111111;
        watermark[2222] <= 18'b111111111111111111;
      end 
      else if((input_valid == 1 || cnt_cycle > 2) && cnt_cycle < 2223) begin
        cnt       <=  cnt + 1;
        cnt_cycle <= cnt / 9;
        wm        <= watermark[cnt_cycle];
      end 
      else begin
        cnt       <= 0;
        cnt_cycle <= 0;
      end 
     
      end
      
      
      
        
 
    

//        Y=0.299*double(R)+0.587*double(G) +0.114*double(B);
//        U=-0.1687*double(R)-0.33163*double(G)+0.5*double(B)+128;
//        V=0.5*double(R)-0.4187*double(G)-0.0813*double(B)+128;

   assign i_imag_Y1[1] = data[576:569] * 306 + data[384:377] * 601 + data[192:185] * 117 ;
   assign i_imag_Y1[2] = data[568:561] * 306 + data[376:369] * 601 + data[184:177] * 117 ;
   assign i_imag_Y1[3] = data[560:553] * 306 + data[368:361] * 601 + data[176:169] * 117 ;
   assign i_imag_Y1[4] = data[552:545] * 306 + data[360:353] * 601 + data[168:161] * 117 ;
   assign i_imag_Y1[5] = data[544:537] * 306 + data[352:345] * 601 + data[160:153] * 117 ;
   assign i_imag_Y1[6] = data[536:529] * 306 + data[344:337] * 601 + data[152:145] * 117 ;
   assign i_imag_Y1[7] = data[528:521] * 306 + data[336:329] * 601 + data[144:137] * 117 ;
   assign i_imag_Y1[8] = data[520:513] * 306 + data[328:321] * 601 + data[136:129] * 117 ;
   assign i_imag_Y2[1] = data[512:505] * 306 + data[320:313] * 601 + data[128:121] * 117 ;
   assign i_imag_Y2[2] = data[504:497] * 306 + data[312:305] * 601 + data[120:113] * 117 ;
   assign i_imag_Y2[3] = data[496:489] * 306 + data[304:297] * 601 + data[112:105] * 117 ;
   assign i_imag_Y2[4] = data[488:481] * 306 + data[296:289] * 601 + data[104:97]  * 117 ;
   assign i_imag_Y2[5] = data[480:473] * 306 + data[288:281] * 601 + data[96:89]   * 117 ;
   assign i_imag_Y2[6] = data[472:465] * 306 + data[280:273] * 601 + data[88:81]   * 117 ;
   assign i_imag_Y2[7] = data[464:457] * 306 + data[272:265] * 601 + data[80:73]   * 117 ;
   assign i_imag_Y2[8] = data[456:449] * 306 + data[264:257] * 601 + data[72:65]   * 117 ;
   assign i_imag_Y3[1] = data[448:441] * 306 + data[256:249] * 601 + data[64:57]   * 117 ;
   assign i_imag_Y3[2] = data[440:433] * 306 + data[248:241] * 601 + data[56:49]   * 117 ;
   assign i_imag_Y3[3] = data[432:425] * 306 + data[240:233] * 601 + data[48:41]   * 117 ;
   assign i_imag_Y3[4] = data[424:417] * 306 + data[232:225] * 601 + data[40:33]   * 117 ;
   assign i_imag_Y3[5] = data[416:409] * 306 + data[224:217] * 601 + data[32:25]   * 117 ;
   assign i_imag_Y3[6] = data[408:401] * 306 + data[216:209] * 601 + data[24:17]   * 117 ;
   assign i_imag_Y3[7] = data[400:393] * 306 + data[208:201] * 601 + data[16:9]    * 117 ;
   assign i_imag_Y3[8] = data[392:385] * 306 + data[200:193] * 601 + data[8:1]     * 117 ;


   assign i_imag_U1[1] = 131072 - data[576:569] * 173 - data[384:377] * 339 + data[192:185] * 512 ;
   assign i_imag_U1[2] = 131072 - data[568:561] * 173 - data[376:369] * 339 + data[184:177] * 512 ;
   assign i_imag_U1[3] = 131072 - data[560:553] * 173 - data[368:361] * 339 + data[176:169] * 512 ;
   assign i_imag_U1[4] = 131072 - data[552:545] * 173 - data[360:353] * 339 + data[168:161] * 512 ;
   assign i_imag_U1[5] = 131072 - data[544:537] * 173 - data[352:345] * 339 + data[160:153] * 512 ;
   assign i_imag_U1[6] = 131072 - data[536:529] * 173 - data[344:337] * 339 + data[152:145] * 512 ;
   assign i_imag_U1[7] = 131072 - data[528:521] * 173 - data[336:329] * 339 + data[144:137] * 512 ;
   assign i_imag_U1[8] = 131072 - data[520:513] * 173 - data[328:321] * 339 + data[136:129] * 512 ;
   assign i_imag_U2[1] = 131072 - data[512:505] * 173 - data[320:313] * 339 + data[128:121] * 512 ;
   assign i_imag_U2[2] = 131072 - data[504:497] * 173 - data[312:305] * 339 + data[120:113] * 512 ;
   assign i_imag_U2[3] = 131072 - data[496:489] * 173 - data[304:297] * 339 + data[112:105] * 512 ;
   assign i_imag_U2[4] = 131072 - data[488:481] * 173 - data[296:289] * 339 + data[104:97]  * 512 ;
   assign i_imag_U2[5] = 131072 - data[480:473] * 173 - data[288:281] * 339 + data[96:89]   * 512 ;
   assign i_imag_U2[6] = 131072 - data[472:465] * 173 - data[280:273] * 339 + data[88:81]   * 512 ;
   assign i_imag_U2[7] = 131072 - data[464:457] * 173 - data[272:265] * 339 + data[80:73]   * 512 ;
   assign i_imag_U2[8] = 131072 - data[456:449] * 173 - data[264:257] * 339 + data[72:65]   * 512 ;
   assign i_imag_U3[1] = 131072 - data[448:441] * 173 - data[256:249] * 339 + data[64:57]   * 512 ;
   assign i_imag_U3[2] = 131072 - data[440:433] * 173 - data[248:241] * 339 + data[56:49]   * 512 ;
   assign i_imag_U3[3] = 131072 - data[432:425] * 173 - data[240:233] * 339 + data[48:41]   * 512 ;
   assign i_imag_U3[4] = 131072 - data[424:417] * 173 - data[232:225] * 339 + data[40:33]   * 512 ;
   assign i_imag_U3[5] = 131072 - data[416:409] * 173 - data[224:217] * 339 + data[32:25]   * 512 ;
   assign i_imag_U3[6] = 131072 - data[408:401] * 173 - data[216:209] * 339 + data[24:17]   * 512 ;
   assign i_imag_U3[7] = 131072 - data[400:393] * 173 - data[208:201] * 339 + data[16:9]    * 512 ;
   assign i_imag_U3[8] = 131072 - data[392:385] * 173 - data[200:193] * 339 + data[8:1]     * 512 ;

   assign i_imag_V1[1] = 131072 + data[576:569] * 512 - data[384:377] * 429 - data[192:185] * 83 ;
   assign i_imag_V1[2] = 131072 + data[568:561] * 512 - data[376:369] * 429 - data[184:177] * 83 ;
   assign i_imag_V1[3] = 131072 + data[560:553] * 512 - data[368:361] * 429 - data[176:169] * 83 ;
   assign i_imag_V1[4] = 131072 + data[552:545] * 512 - data[360:353] * 429 - data[168:161] * 83 ;
   assign i_imag_V1[5] = 131072 + data[544:537] * 512 - data[352:345] * 429 - data[160:153] * 83 ;
   assign i_imag_V1[6] = 131072 + data[536:529] * 512 - data[344:337] * 429 - data[152:145] * 83 ;
   assign i_imag_V1[7] = 131072 + data[528:521] * 512 - data[336:329] * 429 - data[144:137] * 83 ;
   assign i_imag_V1[8] = 131072 + data[520:513] * 512 - data[328:321] * 429 - data[136:129] * 83 ;
   assign i_imag_V2[1] = 131072 + data[512:505] * 512 - data[320:313] * 429 - data[128:121] * 83 ;
   assign i_imag_V2[2] = 131072 + data[504:497] * 512 - data[312:305] * 429 - data[120:113] * 83 ;
   assign i_imag_V2[3] = 131072 + data[496:489] * 512 - data[304:297] * 429 - data[112:105] * 83 ;
   assign i_imag_V2[4] = 131072 + data[488:481] * 512 - data[296:289] * 429 - data[104:97]  * 83 ;
   assign i_imag_V2[5] = 131072 + data[480:473] * 512 - data[288:281] * 429 - data[96:89]   * 83 ;
   assign i_imag_V2[6] = 131072 + data[472:465] * 512 - data[280:273] * 429 - data[88:81]   * 83 ;
   assign i_imag_V2[7] = 131072 + data[464:457] * 512 - data[272:265] * 429 - data[80:73]   * 83 ;
   assign i_imag_V2[8] = 131072 + data[456:449] * 512 - data[264:257] * 429 - data[72:65]   * 83 ;
   assign i_imag_V3[1] = 131072 + data[448:441] * 512 - data[256:249] * 429 - data[64:57]   * 83 ;
   assign i_imag_V3[2] = 131072 + data[440:433] * 512 - data[248:241] * 429 - data[56:49]   * 83 ;
   assign i_imag_V3[3] = 131072 + data[432:425] * 512 - data[240:233] * 429 - data[48:41]   * 83 ;
   assign i_imag_V3[4] = 131072 + data[424:417] * 512 - data[232:225] * 429 - data[40:33]   * 83 ;
   assign i_imag_V3[5] = 131072 + data[416:409] * 512 - data[224:217] * 429 - data[32:25]   * 83 ;
   assign i_imag_V3[6] = 131072 + data[408:401] * 512 - data[216:209] * 429 - data[24:17]   * 83 ;
   assign i_imag_V3[7] = 131072 + data[400:393] * 512 - data[208:201] * 429 - data[16:9]    * 83 ;
   assign i_imag_V3[8] = 131072 + data[392:385] * 512 - data[200:193] * 429 - data[8:1]     * 83 ;


//   R=Y+1.402*(V-128);
//   G=Y-0.34414*(U-128)-0.71414*(V-128);
//   B=Y+1.772*(U-128);
// o_img   8+10
//o_imag_R1
//o_imag_R2
//o_imag_R3
//o_imag_G1
//o_imag_G2
//o_imag_G3
//o_imag_B1
//o_imag_B2
//o_imag_B3

//R1
assign o_imag_R1[1] = o_imag_Y1[1] * 1024 + 1436 * (o_imag_V1[1] - 131072)>0?o_imag_Y1[1] * 1024 + 1436 * (o_imag_V1[1] - 131072):0; 
assign o_imag_R1[2] = o_imag_Y1[2] * 1024 + 1436 * (o_imag_V1[2] - 131072)>0?o_imag_Y1[2] * 1024 + 1436 * (o_imag_V1[2] - 131072):0;
assign o_imag_R1[3] = o_imag_Y1[3] * 1024 + 1436 * (o_imag_V1[3] - 131072)>0?o_imag_Y1[3] * 1024 + 1436 * (o_imag_V1[3] - 131072):0;
assign o_imag_R1[4] = o_imag_Y1[4] * 1024 + 1436 * (o_imag_V1[4] - 131072)>0?o_imag_Y1[4] * 1024 + 1436 * (o_imag_V1[4] - 131072):0;
assign o_imag_R1[5] = o_imag_Y1[5] * 1024 + 1436 * (o_imag_V1[5] - 131072)>0?o_imag_Y1[5] * 1024 + 1436 * (o_imag_V1[5] - 131072):0;
assign o_imag_R1[6] = o_imag_Y1[6] * 1024 + 1436 * (o_imag_V1[6] - 131072)>0?o_imag_Y1[6] * 1024 + 1436 * (o_imag_V1[6] - 131072):0;
assign o_imag_R1[7] = o_imag_Y1[7] * 1024 + 1436 * (o_imag_V1[7] - 131072)>0?o_imag_Y1[7] * 1024 + 1436 * (o_imag_V1[7] - 131072):0;
assign o_imag_R1[8] = o_imag_Y1[8] * 1024 + 1436 * (o_imag_V1[8] - 131072)>0?o_imag_Y1[8] * 1024 + 1436 * (o_imag_V1[8] - 131072):0;
//R2           = o_imag_Y     +      1436 * (= o_imaV_Y   - 131072);      >0?g_Y     +      1436 * (= o_imaV_Y   - 131072);      :0
assign o_imag_R2[1] = o_imag_Y2[1] * 1024 + 1436 * (o_imag_V2[1] - 131072)>0?o_imag_Y2[1] * 1024 + 1436 * (o_imag_V2[1] - 131072):0;
assign o_imag_R2[2] = o_imag_Y2[2] * 1024 + 1436 * (o_imag_V2[2] - 131072)>0?o_imag_Y2[2] * 1024 + 1436 * (o_imag_V2[2] - 131072):0;
assign o_imag_R2[3] = o_imag_Y2[3] * 1024 + 1436 * (o_imag_V2[3] - 131072)>0?o_imag_Y2[3] * 1024 + 1436 * (o_imag_V2[3] - 131072):0;
assign o_imag_R2[4] = o_imag_Y2[4] * 1024 + 1436 * (o_imag_V2[4] - 131072)>0?o_imag_Y2[4] * 1024 + 1436 * (o_imag_V2[4] - 131072):0;
assign o_imag_R2[5] = o_imag_Y2[5] * 1024 + 1436 * (o_imag_V2[5] - 131072)>0?o_imag_Y2[5] * 1024 + 1436 * (o_imag_V2[5] - 131072):0;
assign o_imag_R2[6] = o_imag_Y2[6] * 1024 + 1436 * (o_imag_V2[6] - 131072)>0?o_imag_Y2[6] * 1024 + 1436 * (o_imag_V2[6] - 131072):0;
assign o_imag_R2[7] = o_imag_Y2[7] * 1024 + 1436 * (o_imag_V2[7] - 131072)>0?o_imag_Y2[7] * 1024 + 1436 * (o_imag_V2[7] - 131072):0;
assign o_imag_R2[8] = o_imag_Y2[8] * 1024 + 1436 * (o_imag_V2[8] - 131072)>0?o_imag_Y2[8] * 1024 + 1436 * (o_imag_V2[8] - 131072):0;
 //R3           = o_imag_Y     +      1436 * (= o_imaV_Y   - 131072);     >0?ag_Y     +      1436 * (= o_imaV_Y   - 131072);     :0
assign o_imag_R3[1] = o_imag_Y3[1] * 1024+  1436 * (o_imag_V3[1] - 131072)>0?o_imag_Y3[1] * 1024+  1436 * (o_imag_V3[1] - 131072):0;
assign o_imag_R3[2] = o_imag_Y3[2] * 1024+  1436 * (o_imag_V3[2] - 131072)>0?o_imag_Y3[2] * 1024+  1436 * (o_imag_V3[2] - 131072):0;
assign o_imag_R3[3] = o_imag_Y3[3] * 1024+  1436 * (o_imag_V3[3] - 131072)>0?o_imag_Y3[3] * 1024+  1436 * (o_imag_V3[3] - 131072):0;
assign o_imag_R3[4] = o_imag_Y3[4] * 1024+  1436 * (o_imag_V3[4] - 131072)>0?o_imag_Y3[4] * 1024+  1436 * (o_imag_V3[4] - 131072):0;
assign o_imag_R3[5] = o_imag_Y3[5] * 1024+  1436 * (o_imag_V3[5] - 131072)>0?o_imag_Y3[5] * 1024+  1436 * (o_imag_V3[5] - 131072):0;
assign o_imag_R3[6] = o_imag_Y3[6] * 1024+  1436 * (o_imag_V3[6] - 131072)>0?o_imag_Y3[6] * 1024+  1436 * (o_imag_V3[6] - 131072):0;
assign o_imag_R3[7] = o_imag_Y3[7] * 1024+  1436 * (o_imag_V3[7] - 131072)>0?o_imag_Y3[7] * 1024+  1436 * (o_imag_V3[7] - 131072):0;
assign o_imag_R3[8] = o_imag_Y3[8] * 1024+  1436 * (o_imag_V3[8] - 131072)>0?o_imag_Y3[8] * 1024+  1436 * (o_imag_V3[8] - 131072):0;
//   G=Y-0.34414*(U-128)-0.71414*(V-128);
//G1
assign o_imag_G1[1] = o_imag_Y1[1] * 1024 - 731 * (o_imag_V1[1] - 131072) - 352 * (o_imag_U1[1] - 131072)>0?o_imag_Y1[1] * 1024 - 731 * (o_imag_V1[1] - 131072) - 352 * (o_imag_U1[1] - 131072):0; 
assign o_imag_G1[2] = o_imag_Y1[2] * 1024 - 731 * (o_imag_V1[2] - 131072) - 352 * (o_imag_U1[2] - 131072)>0?o_imag_Y1[2] * 1024 - 731 * (o_imag_V1[2] - 131072) - 352 * (o_imag_U1[2] - 131072):0;
assign o_imag_G1[3] = o_imag_Y1[3] * 1024 - 731 * (o_imag_V1[3] - 131072) - 352 * (o_imag_U1[3] - 131072)>0?o_imag_Y1[3] * 1024 - 731 * (o_imag_V1[3] - 131072) - 352 * (o_imag_U1[3] - 131072):0;
assign o_imag_G1[4] = o_imag_Y1[4] * 1024 - 731 * (o_imag_V1[4] - 131072) - 352 * (o_imag_U1[4] - 131072)>0?o_imag_Y1[4] * 1024 - 731 * (o_imag_V1[4] - 131072) - 352 * (o_imag_U1[4] - 131072):0;
assign o_imag_G1[5] = o_imag_Y1[5] * 1024 - 731 * (o_imag_V1[5] - 131072) - 352 * (o_imag_U1[5] - 131072)>0?o_imag_Y1[5] * 1024 - 731 * (o_imag_V1[5] - 131072) - 352 * (o_imag_U1[5] - 131072):0;
assign o_imag_G1[6] = o_imag_Y1[6] * 1024 - 731 * (o_imag_V1[6] - 131072) - 352 * (o_imag_U1[6] - 131072)>0?o_imag_Y1[6] * 1024 - 731 * (o_imag_V1[6] - 131072) - 352 * (o_imag_U1[6] - 131072):0;
assign o_imag_G1[7] = o_imag_Y1[7] * 1024 - 731 * (o_imag_V1[7] - 131072) - 352 * (o_imag_U1[7] - 131072)>0?o_imag_Y1[7] * 1024 - 731 * (o_imag_V1[7] - 131072) - 352 * (o_imag_U1[7] - 131072):0;
assign o_imag_G1[8] = o_imag_Y1[8] * 1024 - 731 * (o_imag_V1[8] - 131072) - 352 * (o_imag_U1[8] - 131072)>0?o_imag_Y1[8] * 1024 - 731 * (o_imag_V1[8] - 131072) - 352 * (o_imag_U1[8] - 131072):0;
 //G2   G       = o_imag_Y     +    - 731 * (= o_imaV_Y   - 131072) - 352 * (= o_imaU_Y   - 131072);     >0?ag_Y     +    - 731 * (= o_imaV_Y   - 131072) - 352 * (= o_imaU_Y   - 131072);     :0
assign o_imag_G2[1] = o_imag_Y2[1] * 1024 - 731 * (o_imag_V2[1] - 131072) - 352 * (o_imag_U2[1] - 131072)>0?o_imag_Y2[1] * 1024 - 731 * (o_imag_V2[1] - 131072) - 352 * (o_imag_U2[1] - 131072):0;
assign o_imag_G2[2] = o_imag_Y2[2] * 1024 - 731 * (o_imag_V2[2] - 131072) - 352 * (o_imag_U2[2] - 131072)>0?o_imag_Y2[2] * 1024 - 731 * (o_imag_V2[2] - 131072) - 352 * (o_imag_U2[2] - 131072):0;
assign o_imag_G2[3] = o_imag_Y2[3] * 1024 - 731 * (o_imag_V2[3] - 131072) - 352 * (o_imag_U2[3] - 131072)>0?o_imag_Y2[3] * 1024 - 731 * (o_imag_V2[3] - 131072) - 352 * (o_imag_U2[3] - 131072):0;
assign o_imag_G2[4] = o_imag_Y2[4] * 1024 - 731 * (o_imag_V2[4] - 131072) - 352 * (o_imag_U2[4] - 131072)>0?o_imag_Y2[4] * 1024 - 731 * (o_imag_V2[4] - 131072) - 352 * (o_imag_U2[4] - 131072):0;
assign o_imag_G2[5] = o_imag_Y2[5] * 1024 - 731 * (o_imag_V2[5] - 131072) - 352 * (o_imag_U2[5] - 131072)>0?o_imag_Y2[5] * 1024 - 731 * (o_imag_V2[5] - 131072) - 352 * (o_imag_U2[5] - 131072):0;
assign o_imag_G2[6] = o_imag_Y2[6] * 1024 - 731 * (o_imag_V2[6] - 131072) - 352 * (o_imag_U2[6] - 131072)>0?o_imag_Y2[6] * 1024 - 731 * (o_imag_V2[6] - 131072) - 352 * (o_imag_U2[6] - 131072):0;
assign o_imag_G2[7] = o_imag_Y2[7] * 1024 - 731 * (o_imag_V2[7] - 131072) - 352 * (o_imag_U2[7] - 131072)>0?o_imag_Y2[7] * 1024 - 731 * (o_imag_V2[7] - 131072) - 352 * (o_imag_U2[7] - 131072):0;
assign o_imag_G2[8] = o_imag_Y2[8] * 1024 - 731 * (o_imag_V2[8] - 131072) - 352 * (o_imag_U2[8] - 131072)>0?o_imag_Y2[8] * 1024 - 731 * (o_imag_V2[8] - 131072) - 352 * (o_imag_U2[8] - 131072):0;
//G3   G       = o_imag_Y     +    - 731 * (= o_imaV_Y   - 131072) - 352 * (= o_imaU_Y   - 131072);      >0?g_Y     +    - 731 * (= o_imaV_Y   - 131072) - 352 * (= o_imaU_Y   - 131072);      :0
assign o_imag_G3[1] = o_imag_Y3[1] * 1024 - 731 * (o_imag_V3[1] - 131072) - 352 * (o_imag_U3[1] - 131072)>0?o_imag_Y3[1] * 1024 - 731 * (o_imag_V3[1] - 131072) - 352 * (o_imag_U3[1] - 131072):0;
assign o_imag_G3[2] = o_imag_Y3[2] * 1024 - 731 * (o_imag_V3[2] - 131072) - 352 * (o_imag_U3[2] - 131072)>0?o_imag_Y3[2] * 1024 - 731 * (o_imag_V3[2] - 131072) - 352 * (o_imag_U3[2] - 131072):0;
assign o_imag_G3[3] = o_imag_Y3[3] * 1024 - 731 * (o_imag_V3[3] - 131072) - 352 * (o_imag_U3[3] - 131072)>0?o_imag_Y3[3] * 1024 - 731 * (o_imag_V3[3] - 131072) - 352 * (o_imag_U3[3] - 131072):0;
assign o_imag_G3[4] = o_imag_Y3[4] * 1024 - 731 * (o_imag_V3[4] - 131072) - 352 * (o_imag_U3[4] - 131072)>0?o_imag_Y3[4] * 1024 - 731 * (o_imag_V3[4] - 131072) - 352 * (o_imag_U3[4] - 131072):0;
assign o_imag_G3[5] = o_imag_Y3[5] * 1024 - 731 * (o_imag_V3[5] - 131072) - 352 * (o_imag_U3[5] - 131072)>0?o_imag_Y3[5] * 1024 - 731 * (o_imag_V3[5] - 131072) - 352 * (o_imag_U3[5] - 131072):0;
assign o_imag_G3[6] = o_imag_Y3[6] * 1024 - 731 * (o_imag_V3[6] - 131072) - 352 * (o_imag_U3[6] - 131072)>0?o_imag_Y3[6] * 1024 - 731 * (o_imag_V3[6] - 131072) - 352 * (o_imag_U3[6] - 131072):0;
assign o_imag_G3[7] = o_imag_Y3[7] * 1024 - 731 * (o_imag_V3[7] - 131072) - 352 * (o_imag_U3[7] - 131072)>0?o_imag_Y3[7] * 1024 - 731 * (o_imag_V3[7] - 131072) - 352 * (o_imag_U3[7] - 131072):0;
assign o_imag_G3[8] = o_imag_Y3[8] * 1024 - 731 * (o_imag_V3[8] - 131072) - 352 * (o_imag_U3[8] - 131072)>0?o_imag_Y3[8] * 1024 - 731 * (o_imag_V3[8] - 131072) - 352 * (o_imag_U3[8] - 131072):0;
//   B=Y+1.772*(U-128);                                                               
//R1
assign o_imag_B1[1] = o_imag_Y1[1] * 1024 + 1814 * (o_imag_U1[1] - 131072)>0?o_imag_Y1[1] * 1024 + 1814 * (o_imag_U1[1] - 131072):0; 
assign o_imag_B1[2] = o_imag_Y1[2] * 1024 + 1814 * (o_imag_U1[2] - 131072)>0?o_imag_Y1[2] * 1024 + 1814 * (o_imag_U1[2] - 131072):0;
assign o_imag_B1[3] = o_imag_Y1[3] * 1024 + 1814 * (o_imag_U1[3] - 131072)>0?o_imag_Y1[3] * 1024 + 1814 * (o_imag_U1[3] - 131072):0;
assign o_imag_B1[4] = o_imag_Y1[4] * 1024 + 1814 * (o_imag_U1[4] - 131072)>0?o_imag_Y1[4] * 1024 + 1814 * (o_imag_U1[4] - 131072):0;
assign o_imag_B1[5] = o_imag_Y1[5] * 1024 + 1814 * (o_imag_U1[5] - 131072)>0?o_imag_Y1[5] * 1024 + 1814 * (o_imag_U1[5] - 131072):0;
assign o_imag_B1[6] = o_imag_Y1[6] * 1024 + 1814 * (o_imag_U1[6] - 131072)>0?o_imag_Y1[6] * 1024 + 1814 * (o_imag_U1[6] - 131072):0;
assign o_imag_B1[7] = o_imag_Y1[7] * 1024 + 1814 * (o_imag_U1[7] - 131072)>0?o_imag_Y1[7] * 1024 + 1814 * (o_imag_U1[7] - 131072):0;
assign o_imag_B1[8] = o_imag_Y1[8] * 1024 + 1814 * (o_imag_U1[8] - 131072)>0?o_imag_Y1[8] * 1024 + 1814 * (o_imag_U1[8] - 131072):0;
//R2   B       = o_imag_Y     +      1814 * (= o_imaU_Y   - 131072);      >0?g_Y     +      1814 * (= o_imaU_Y   - 131072);      :0
assign o_imag_B2[1] = o_imag_Y2[1] * 1024 + 1814 * (o_imag_U2[1] - 131072)>0?o_imag_Y2[1] * 1024 + 1814 * (o_imag_U2[1] - 131072):0;
assign o_imag_B2[2] = o_imag_Y2[2] * 1024 + 1814 * (o_imag_U2[2] - 131072)>0?o_imag_Y2[2] * 1024 + 1814 * (o_imag_U2[2] - 131072):0;
assign o_imag_B2[3] = o_imag_Y2[3] * 1024 + 1814 * (o_imag_U2[3] - 131072)>0?o_imag_Y2[3] * 1024 + 1814 * (o_imag_U2[3] - 131072):0;
assign o_imag_B2[4] = o_imag_Y2[4] * 1024 + 1814 * (o_imag_U2[4] - 131072)>0?o_imag_Y2[4] * 1024 + 1814 * (o_imag_U2[4] - 131072):0;
assign o_imag_B2[5] = o_imag_Y2[5] * 1024 + 1814 * (o_imag_U2[5] - 131072)>0?o_imag_Y2[5] * 1024 + 1814 * (o_imag_U2[5] - 131072):0;
assign o_imag_B2[6] = o_imag_Y2[6] * 1024 + 1814 * (o_imag_U2[6] - 131072)>0?o_imag_Y2[6] * 1024 + 1814 * (o_imag_U2[6] - 131072):0;
assign o_imag_B2[7] = o_imag_Y2[7] * 1024 + 1814 * (o_imag_U2[7] - 131072)>0?o_imag_Y2[7] * 1024 + 1814 * (o_imag_U2[7] - 131072):0;
assign o_imag_B2[8] = o_imag_Y2[8] * 1024 + 1814 * (o_imag_U2[8] - 131072)>0?o_imag_Y2[8] * 1024 + 1814 * (o_imag_U2[8] - 131072):0;
 //R3   B       = o_imag_Y     +      1814 * (= o_imaU_Y   - 131072);     >0?ag_Y     +      1814 * (= o_imaU_Y   - 131072);     :0
assign o_imag_B3[1] = o_imag_Y3[1] * 1024+  1814 * (o_imag_U3[1] - 131072)>0?o_imag_Y3[1] * 1024+  1814 * (o_imag_U3[1] - 131072):0;
assign o_imag_B3[2] = o_imag_Y3[2] * 1024+  1814 * (o_imag_U3[2] - 131072)>0?o_imag_Y3[2] * 1024+  1814 * (o_imag_U3[2] - 131072):0;
assign o_imag_B3[3] = o_imag_Y3[3] * 1024+  1814 * (o_imag_U3[3] - 131072)>0?o_imag_Y3[3] * 1024+  1814 * (o_imag_U3[3] - 131072):0;
assign o_imag_B3[4] = o_imag_Y3[4] * 1024+  1814 * (o_imag_U3[4] - 131072)>0?o_imag_Y3[4] * 1024+  1814 * (o_imag_U3[4] - 131072):0;
assign o_imag_B3[5] = o_imag_Y3[5] * 1024+  1814 * (o_imag_U3[5] - 131072)>0?o_imag_Y3[5] * 1024+  1814 * (o_imag_U3[5] - 131072):0;
assign o_imag_B3[6] = o_imag_Y3[6] * 1024+  1814 * (o_imag_U3[6] - 131072)>0?o_imag_Y3[6] * 1024+  1814 * (o_imag_U3[6] - 131072):0;
assign o_imag_B3[7] = o_imag_Y3[7] * 1024+  1814 * (o_imag_U3[7] - 131072)>0?o_imag_Y3[7] * 1024+  1814 * (o_imag_U3[7] - 131072):0;
assign o_imag_B3[8] = o_imag_Y3[8] * 1024+  1814 * (o_imag_U3[8] - 131072)>0?o_imag_Y3[8] * 1024+  1814 * (o_imag_U3[8] - 131072):0;

assign o_data = { o_imag_R1_f[1],o_imag_R1_f[2],o_imag_R1_f[3],o_imag_R1_f[4],o_imag_R1_f[5],o_imag_R1_f[6],o_imag_R1_f[7],o_imag_R1_f[8],
                  o_imag_R2_f[1],o_imag_R2_f[2],o_imag_R2_f[3],o_imag_R2_f[4],o_imag_R2_f[5],o_imag_R2_f[6],o_imag_R2_f[7],o_imag_R2_f[8],
                  o_imag_R3_f[1],o_imag_R3_f[2],o_imag_R3_f[3],o_imag_R3_f[4],o_imag_R3_f[5],o_imag_R3_f[6],o_imag_R3_f[7],o_imag_R3_f[8],   
                  o_imag_G1_f[1],o_imag_G1_f[2],o_imag_G1_f[3],o_imag_G1_f[4],o_imag_G1_f[5],o_imag_G1_f[6],o_imag_G1_f[7],o_imag_G1_f[8],   
                  o_imag_G2_f[1],o_imag_G2_f[2],o_imag_G2_f[3],o_imag_G2_f[4],o_imag_G2_f[5],o_imag_G2_f[6],o_imag_G2_f[7],o_imag_G2_f[8],   
                  o_imag_G3_f[1],o_imag_G3_f[2],o_imag_G3_f[3],o_imag_G3_f[4],o_imag_G3_f[5],o_imag_G3_f[6],o_imag_G3_f[7],o_imag_G3_f[8],      
                  o_imag_B1_f[1],o_imag_B1_f[2],o_imag_B1_f[3],o_imag_B1_f[4],o_imag_B1_f[5],o_imag_B1_f[6],o_imag_B1_f[7],o_imag_B1_f[8], 
                  o_imag_B2_f[1],o_imag_B2_f[2],o_imag_B2_f[3],o_imag_B2_f[4],o_imag_B2_f[5],o_imag_B2_f[6],o_imag_B2_f[7],o_imag_B2_f[8], 
                  o_imag_B3_f[1],o_imag_B3_f[2],o_imag_B3_f[3],o_imag_B3_f[4],o_imag_B3_f[5],o_imag_B3_f[6],o_imag_B3_f[7],o_imag_B3_f[8]
                 };


     wmins_4 CAL_Y1(

               .clk   (clk),
               .rst   (rst),

               .image_1( i_imag_Y1[1]),//1+8+0  {signal,0-255}
               .image_2( i_imag_Y1[2]),
               .image_3( i_imag_Y1[3]),
               .image_4( i_imag_Y1[4]),
               .image_5( i_imag_Y1[5]),
               .image_6( i_imag_Y1[6]),
               .image_7( i_imag_Y1[7]),
               .image_8( i_imag_Y1[8]),

               .ins_M  (/*wm[18:15]*/4'b1011),


               .image_ins_1(o_imag_Y1[1][18:1]),
               .image_ins_2(o_imag_Y1[2][18:1]),
               .image_ins_3(o_imag_Y1[3][18:1]),
               .image_ins_4(o_imag_Y1[4][18:1]),
               .image_ins_5(o_imag_Y1[5][18:1]),
               .image_ins_6(o_imag_Y1[6][18:1]),
               .image_ins_7(o_imag_Y1[7][18:1]),
               .image_ins_8(o_imag_Y1[8][18:1]),

               .ins_mode  (1'b0         ),
               .input_valid(input_valid),
               .output_valid()



                   );

      wmins_4 CAL_Y2(

               .clk   (clk),
               .rst   (rst),

               .image_1( i_imag_Y2[1]),//1+8+0  {signal,0-255}
               .image_2( i_imag_Y2[2]),
               .image_3( i_imag_Y2[3]),
               .image_4( i_imag_Y2[4]),
               .image_5( i_imag_Y2[5]),
               .image_6( i_imag_Y2[6]),
               .image_7( i_imag_Y2[7]),
               .image_8( i_imag_Y2[8]),

               .ins_M  (wm[14:11]),


               .image_ins_1(o_imag_Y2[1][18:1]),
               .image_ins_2(o_imag_Y2[2][18:1]),
               .image_ins_3(o_imag_Y2[3][18:1]),
               .image_ins_4(o_imag_Y2[4][18:1]),
               .image_ins_5(o_imag_Y2[5][18:1]),
               .image_ins_6(o_imag_Y2[6][18:1]),
               .image_ins_7(o_imag_Y2[7][18:1]),
               .image_ins_8(o_imag_Y2[8][18:1]),

               .ins_mode  (1'b0         ),
               .input_valid(input_valid),
               .output_valid()



                   );


            wmins_4 CAL_Y3(

               .clk   (clk),
               .rst   (rst),

               .image_1( i_imag_Y3[1]),//1+8+0  {signal,0-255}
               .image_2( i_imag_Y3[2]),
               .image_3( i_imag_Y3[3]),
               .image_4( i_imag_Y3[4]),
               .image_5( i_imag_Y3[5]),
               .image_6( i_imag_Y3[6]),
               .image_7( i_imag_Y3[7]),
               .image_8( i_imag_Y3[8]),

               .ins_M  (wm[10:7]),


               .image_ins_1(o_imag_Y3[1][18:1]),
               .image_ins_2(o_imag_Y3[2][18:1]),
               .image_ins_3(o_imag_Y3[3][18:1]),
               .image_ins_4(o_imag_Y3[4][18:1]),
               .image_ins_5(o_imag_Y3[5][18:1]),
               .image_ins_6(o_imag_Y3[6][18:1]),
               .image_ins_7(o_imag_Y3[7][18:1]),
               .image_ins_8(o_imag_Y3[8][18:1]),

               .ins_mode  (1'b0         ),
               .input_valid(input_valid),
               .output_valid()



                   );

             wmins_4 CAL_U1(

               .clk   (clk),
               .rst   (rst),

               .image_1( i_imag_U1[1]),//1+8+0  {signal,0-255}
               .image_2( i_imag_U1[2]),
               .image_3( i_imag_U1[3]),
               .image_4( i_imag_U1[4]),
               .image_5( i_imag_U1[5]),
               .image_6( i_imag_U1[6]),
               .image_7( i_imag_U1[7]),
               .image_8( i_imag_U1[8]),

               .ins_M  ({4'b0001}),
//wm[6]

               .image_ins_1(o_imag_U1[1][18:1]),
               .image_ins_2(o_imag_U1[2][18:1]),
               .image_ins_3(o_imag_U1[3][18:1]),
               .image_ins_4(o_imag_U1[4][18:1]),
               .image_ins_5(o_imag_U1[5][18:1]),
               .image_ins_6(o_imag_U1[6][18:1]),
               .image_ins_7(o_imag_U1[7][18:1]),
               .image_ins_8(o_imag_U1[8][18:1]),

               .ins_mode  (1'b1         ),
               .input_valid(input_valid),
               .output_valid()



                   );

             wmins_4 CAL_U2(

               .clk   (clk),
               .rst   (rst),

               .image_1( i_imag_U2[1]),//1+8+0  {signal,0-255}
               .image_2( i_imag_U2[2]),
               .image_3( i_imag_U2[3]),
               .image_4( i_imag_U2[4]),
               .image_5( i_imag_U2[5]),
               .image_6( i_imag_U2[6]),
               .image_7( i_imag_U2[7]),
               .image_8( i_imag_U2[8]),

               .ins_M  ({3'b000,wm[5]}),


               .image_ins_1(o_imag_U2[1][18:1]),
               .image_ins_2(o_imag_U2[2][18:1]),
               .image_ins_3(o_imag_U2[3][18:1]),
               .image_ins_4(o_imag_U2[4][18:1]),
               .image_ins_5(o_imag_U2[5][18:1]),
               .image_ins_6(o_imag_U2[6][18:1]),
               .image_ins_7(o_imag_U2[7][18:1]),
               .image_ins_8(o_imag_U2[8][18:1]),

               .ins_mode  (1'b1         ),
               .input_valid(input_valid),
               .output_valid()



                   );

             wmins_4 CAL_U3(

               .clk   (clk),
               .rst   (rst),

               .image_1( i_imag_U3[1]),//1+8+0  {signal,0-255}
               .image_2( i_imag_U3[2]),
               .image_3( i_imag_U3[3]),
               .image_4( i_imag_U3[4]),
               .image_5( i_imag_U3[5]),
               .image_6( i_imag_U3[6]),
               .image_7( i_imag_U3[7]),
               .image_8( i_imag_U3[8]),

               .ins_M  ({3'b000,wm[4]}),


               .image_ins_1(o_imag_U3[1][18:1]),
               .image_ins_2(o_imag_U3[2][18:1]),
               .image_ins_3(o_imag_U3[3][18:1]),
               .image_ins_4(o_imag_U3[4][18:1]),
               .image_ins_5(o_imag_U3[5][18:1]),
               .image_ins_6(o_imag_U3[6][18:1]),
               .image_ins_7(o_imag_U3[7][18:1]),
               .image_ins_8(o_imag_U3[8][18:1]),

               .ins_mode  (1'b1         ),
               .input_valid(input_valid),
               .output_valid()



                   );

             wmins_4 CAL_V1(

               .clk   (clk),
               .rst   (rst),

               .image_1( i_imag_V1[1]),//1+8+0  {signal,0-255}
               .image_2( i_imag_V1[2]),
               .image_3( i_imag_V1[3]),
               .image_4( i_imag_V1[4]),
               .image_5( i_imag_V1[5]),
               .image_6( i_imag_V1[6]),
               .image_7( i_imag_V1[7]),
               .image_8( i_imag_V1[8]),

               .ins_M  ({4'b0001}),


               .image_ins_1(o_imag_V1[1][18:1]),
               .image_ins_2(o_imag_V1[2][18:1]),
               .image_ins_3(o_imag_V1[3][18:1]),
               .image_ins_4(o_imag_V1[4][18:1]),
               .image_ins_5(o_imag_V1[5][18:1]),
               .image_ins_6(o_imag_V1[6][18:1]),
               .image_ins_7(o_imag_V1[7][18:1]),
               .image_ins_8(o_imag_V1[8][18:1]),

               .ins_mode  (1'b1         ),
               .input_valid(input_valid),
               .output_valid()



                   );

             wmins_4 CAL_V2(

               .clk   (clk),
               .rst   (rst),

               .image_1( i_imag_V2[1]),//1+8+0  {signal,0-255}
               .image_2( i_imag_V2[2]),
               .image_3( i_imag_V2[3]),
               .image_4( i_imag_V2[4]),
               .image_5( i_imag_V2[5]),
               .image_6( i_imag_V2[6]),
               .image_7( i_imag_V2[7]),
               .image_8( i_imag_V2[8]),

               .ins_M  ({3'b000,wm[2]}),


               .image_ins_1(o_imag_V2[1][18:1]),
               .image_ins_2(o_imag_V2[2][18:1]),
               .image_ins_3(o_imag_V2[3][18:1]),
               .image_ins_4(o_imag_V2[4][18:1]),
               .image_ins_5(o_imag_V2[5][18:1]),
               .image_ins_6(o_imag_V2[6][18:1]),
               .image_ins_7(o_imag_V2[7][18:1]),
               .image_ins_8(o_imag_V2[8][18:1]),

               .ins_mode  (1'b1         ),
               .input_valid(input_valid),
               .output_valid()



                   );

             wmins_4 CAL_V3(

               .clk   (clk),
               .rst   (rst),

               .image_1( i_imag_V3[1]),//1+8+0  {signal,0-255}
               .image_2( i_imag_V3[2]),
               .image_3( i_imag_V3[3]),
               .image_4( i_imag_V3[4]),
               .image_5( i_imag_V3[5]),
               .image_6( i_imag_V3[6]),
               .image_7( i_imag_V3[7]),
               .image_8( i_imag_V3[8]),

               .ins_M  ({3'b000,wm[1]}),


               .image_ins_1(o_imag_V3[1][18:1]),
               .image_ins_2(o_imag_V3[2][18:1]),
               .image_ins_3(o_imag_V3[3][18:1]),
               .image_ins_4(o_imag_V3[4][18:1]),
               .image_ins_5(o_imag_V3[5][18:1]),
               .image_ins_6(o_imag_V3[6][18:1]),
               .image_ins_7(o_imag_V3[7][18:1]),
               .image_ins_8(o_imag_V3[8][18:1]),

               .ins_mode  (1'b1         ),
               .input_valid(input_valid),
               .output_valid()



                   );
                   
   watermark_dataset inst(
                            .clk   (clk) ,
                            .valid (input_valid) ,
                            .rst   (rst) ,
                            .o_data(data)
                            );

endmodule
