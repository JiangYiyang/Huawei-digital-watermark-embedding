`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/08/17 23:58:24
// Design Name: 
// Module Name: cossin_24
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module cossin_24(
    
    input wire signed [24:1] rad,
    output  wire signed [24:1] cos,
    output  wire signed [24:1] sin
        );
    wire [1:0] sig ;
    wire signed [24:1] rad_abs;
    wire signed [24:1] rad_abs_90;
    reg signed [24:1] cos_tmp;
    reg signed [24:1] sin_tmp;
    
    assign sig = {rad[24],rad_abs[24:13] > 805};
    assign rad_abs = sig[1] ? - rad : rad ;
    assign rad_abs_90 = sig[0] ? 24'd6588397- rad_abs : rad_abs; 
    assign cos = sig[0] ? - cos_tmp : cos_tmp  ;
    assign sin = sig[1] ? - sin_tmp : sin_tmp  ;
    always @(*) begin
      case(rad_abs_90[24:13])
      12'd0: begin cos_tmp = 24'b001111111111111111101011 ; sin_tmp = 24'b000000000011001101111001 ; end 
      12'd1: begin cos_tmp = 24'b001111111111111111101011 ; sin_tmp = 24'b000000000011001101111001 ; end 
      12'd2: begin cos_tmp = 24'b001111111111111110101101 ; sin_tmp = 24'b000000000110011011110001 ; end 
      12'd3: begin cos_tmp = 24'b001111111111111101000110 ; sin_tmp = 24'b000000001001101001101010 ; end 
      12'd4: begin cos_tmp = 24'b001111111111111101000110 ; sin_tmp = 24'b000000001001101001101010 ; end 
      12'd5: begin cos_tmp = 24'b001111111111111010110101 ; sin_tmp = 24'b000000001100110111100010 ; end 
      12'd6: begin cos_tmp = 24'b001111111111110111111011 ; sin_tmp = 24'b000000010000000101011001 ; end 
      12'd7: begin cos_tmp = 24'b001111111111110111111011 ; sin_tmp = 24'b000000010000000101011001 ; end 
      12'd8: begin cos_tmp = 24'b001111111111110100010111 ; sin_tmp = 24'b000000010011010011010000 ; end 
      12'd9: begin cos_tmp = 24'b001111111111110100010111 ; sin_tmp = 24'b000000010011010011010000 ; end 
      12'd10: begin cos_tmp = 24'b001111111111110000001010 ; sin_tmp = 24'b000000010110100001000110 ; end 
      12'd11: begin cos_tmp = 24'b001111111111101011010011 ; sin_tmp = 24'b000000011001101110111011 ; end 
      12'd12: begin cos_tmp = 24'b001111111111101011010011 ; sin_tmp = 24'b000000011001101110111011 ; end 
      12'd13: begin cos_tmp = 24'b001111111111100101110100 ; sin_tmp = 24'b000000011100111100101111 ; end 
      12'd14: begin cos_tmp = 24'b001111111111011111101010 ; sin_tmp = 24'b000000100000001010100010 ; end 
      12'd15: begin cos_tmp = 24'b001111111111011111101010 ; sin_tmp = 24'b000000100000001010100010 ; end 
      12'd16: begin cos_tmp = 24'b001111111111011000111000 ; sin_tmp = 24'b000000100011011000010100 ; end 
      12'd17: begin cos_tmp = 24'b001111111111011000111000 ; sin_tmp = 24'b000000100011011000010100 ; end 
      12'd18: begin cos_tmp = 24'b001111111111010001011100 ; sin_tmp = 24'b000000100110100110000100 ; end 
      12'd19: begin cos_tmp = 24'b001111111111001001010111 ; sin_tmp = 24'b000000101001110011110011 ; end 
      12'd20: begin cos_tmp = 24'b001111111111001001010111 ; sin_tmp = 24'b000000101001110011110011 ; end 
      12'd21: begin cos_tmp = 24'b001111111111000000101000 ; sin_tmp = 24'b000000101101000001100000 ; end 
      12'd22: begin cos_tmp = 24'b001111111111000000101000 ; sin_tmp = 24'b000000101101000001100000 ; end 
      12'd23: begin cos_tmp = 24'b001111111110110111010000 ; sin_tmp = 24'b000000110000001111001011 ; end 
      12'd24: begin cos_tmp = 24'b001111111110101101001110 ; sin_tmp = 24'b000000110011011100110100 ; end 
      12'd25: begin cos_tmp = 24'b001111111110101101001110 ; sin_tmp = 24'b000000110011011100110100 ; end 
      12'd26: begin cos_tmp = 24'b001111111110100010100100 ; sin_tmp = 24'b000000110110101010011011 ; end 
      12'd27: begin cos_tmp = 24'b001111111110010111010000 ; sin_tmp = 24'b000000111001111000000000 ; end 
      12'd28: begin cos_tmp = 24'b001111111110010111010000 ; sin_tmp = 24'b000000111001111000000000 ; end 
      12'd29: begin cos_tmp = 24'b001111111110001011010010 ; sin_tmp = 24'b000000111101000101100010 ; end 
      12'd30: begin cos_tmp = 24'b001111111110001011010010 ; sin_tmp = 24'b000000111101000101100010 ; end 
      12'd31: begin cos_tmp = 24'b001111111101111110101011 ; sin_tmp = 24'b000001000000010011000011 ; end 
      12'd32: begin cos_tmp = 24'b001111111101110001011011 ; sin_tmp = 24'b000001000011100000100000 ; end 
      12'd33: begin cos_tmp = 24'b001111111101110001011011 ; sin_tmp = 24'b000001000011100000100000 ; end 
      12'd34: begin cos_tmp = 24'b001111111101100011100010 ; sin_tmp = 24'b000001000110101101111011 ; end 
      12'd35: begin cos_tmp = 24'b001111111101010100111111 ; sin_tmp = 24'b000001001001111011010011 ; end 
      12'd36: begin cos_tmp = 24'b001111111101010100111111 ; sin_tmp = 24'b000001001001111011010011 ; end 
      12'd37: begin cos_tmp = 24'b001111111101000101110100 ; sin_tmp = 24'b000001001101001000101000 ; end 
      12'd38: begin cos_tmp = 24'b001111111101000101110100 ; sin_tmp = 24'b000001001101001000101000 ; end 
      12'd39: begin cos_tmp = 24'b001111111100110101111110 ; sin_tmp = 24'b000001010000010101111001 ; end 
      12'd40: begin cos_tmp = 24'b001111111100100101100000 ; sin_tmp = 24'b000001010011100011001000 ; end 
      12'd41: begin cos_tmp = 24'b001111111100100101100000 ; sin_tmp = 24'b000001010011100011001000 ; end 
      12'd42: begin cos_tmp = 24'b001111111100010100011000 ; sin_tmp = 24'b000001010110110000010011 ; end 
      12'd43: begin cos_tmp = 24'b001111111100000010100111 ; sin_tmp = 24'b000001011001111101011011 ; end 
      12'd44: begin cos_tmp = 24'b001111111100000010100111 ; sin_tmp = 24'b000001011001111101011011 ; end 
      12'd45: begin cos_tmp = 24'b001111111011110000001101 ; sin_tmp = 24'b000001011101001010011111 ; end 
      12'd46: begin cos_tmp = 24'b001111111011110000001101 ; sin_tmp = 24'b000001011101001010011111 ; end 
      12'd47: begin cos_tmp = 24'b001111111011011101001010 ; sin_tmp = 24'b000001100000010111011111 ; end 
      12'd48: begin cos_tmp = 24'b001111111011001001011101 ; sin_tmp = 24'b000001100011100100011011 ; end 
      12'd49: begin cos_tmp = 24'b001111111011001001011101 ; sin_tmp = 24'b000001100011100100011011 ; end 
      12'd50: begin cos_tmp = 24'b001111111010110101000111 ; sin_tmp = 24'b000001100110110001010100 ; end 
      12'd51: begin cos_tmp = 24'b001111111010100000001000 ; sin_tmp = 24'b000001101001111110001000 ; end 
      12'd52: begin cos_tmp = 24'b001111111010100000001000 ; sin_tmp = 24'b000001101001111110001000 ; end 
      12'd53: begin cos_tmp = 24'b001111111010001010100000 ; sin_tmp = 24'b000001101101001010111000 ; end 
      12'd54: begin cos_tmp = 24'b001111111010001010100000 ; sin_tmp = 24'b000001101101001010111000 ; end 
      12'd55: begin cos_tmp = 24'b001111111001110100001110 ; sin_tmp = 24'b000001110000010111100011 ; end 
      12'd56: begin cos_tmp = 24'b001111111001011101010100 ; sin_tmp = 24'b000001110011100100001010 ; end 
      12'd57: begin cos_tmp = 24'b001111111001011101010100 ; sin_tmp = 24'b000001110011100100001010 ; end 
      12'd58: begin cos_tmp = 24'b001111111001000101110000 ; sin_tmp = 24'b000001110110110000101100 ; end 
      12'd59: begin cos_tmp = 24'b001111111001000101110000 ; sin_tmp = 24'b000001110110110000101100 ; end 
      12'd60: begin cos_tmp = 24'b001111111000101101100011 ; sin_tmp = 24'b000001111001111101001010 ; end 
      12'd61: begin cos_tmp = 24'b001111111000010100101110 ; sin_tmp = 24'b000001111101001001100010 ; end 
      12'd62: begin cos_tmp = 24'b001111111000010100101110 ; sin_tmp = 24'b000001111101001001100010 ; end 
      12'd63: begin cos_tmp = 24'b001111110111111011001111 ; sin_tmp = 24'b000010000000010101110110 ; end 
      12'd64: begin cos_tmp = 24'b001111110111100001000111 ; sin_tmp = 24'b000010000011100010000100 ; end 
      12'd65: begin cos_tmp = 24'b001111110111100001000111 ; sin_tmp = 24'b000010000011100010000100 ; end 
      12'd66: begin cos_tmp = 24'b001111110111000110010110 ; sin_tmp = 24'b000010000110101110001101 ; end 
      12'd67: begin cos_tmp = 24'b001111110111000110010110 ; sin_tmp = 24'b000010000110101110001101 ; end 
      12'd68: begin cos_tmp = 24'b001111110110101010111011 ; sin_tmp = 24'b000010001001111010010000 ; end 
      12'd69: begin cos_tmp = 24'b001111110110001110111000 ; sin_tmp = 24'b000010001101000110001110 ; end 
      12'd70: begin cos_tmp = 24'b001111110110001110111000 ; sin_tmp = 24'b000010001101000110001110 ; end 
      12'd71: begin cos_tmp = 24'b001111110101110010001100 ; sin_tmp = 24'b000010010000010010000111 ; end 
      12'd72: begin cos_tmp = 24'b001111110101010100110111 ; sin_tmp = 24'b000010010011011101111001 ; end 
      12'd73: begin cos_tmp = 24'b001111110101010100110111 ; sin_tmp = 24'b000010010011011101111001 ; end 
      12'd74: begin cos_tmp = 24'b001111110100110110111001 ; sin_tmp = 24'b000010010110101001100101 ; end 
      12'd75: begin cos_tmp = 24'b001111110100110110111001 ; sin_tmp = 24'b000010010110101001100101 ; end 
      12'd76: begin cos_tmp = 24'b001111110100011000010010 ; sin_tmp = 24'b000010011001110101001100 ; end 
      12'd77: begin cos_tmp = 24'b001111110011111001000010 ; sin_tmp = 24'b000010011101000000101100 ; end 
      12'd78: begin cos_tmp = 24'b001111110011111001000010 ; sin_tmp = 24'b000010011101000000101100 ; end 
      12'd79: begin cos_tmp = 24'b001111110011011001001001 ; sin_tmp = 24'b000010100000001100000110 ; end 
      12'd80: begin cos_tmp = 24'b001111110010111000100111 ; sin_tmp = 24'b000010100011010111011001 ; end 
      12'd81: begin cos_tmp = 24'b001111110010111000100111 ; sin_tmp = 24'b000010100011010111011001 ; end 
      12'd82: begin cos_tmp = 24'b001111110010010111011101 ; sin_tmp = 24'b000010100110100010100110 ; end 
      12'd83: begin cos_tmp = 24'b001111110010010111011101 ; sin_tmp = 24'b000010100110100010100110 ; end 
      12'd84: begin cos_tmp = 24'b001111110001110101101001 ; sin_tmp = 24'b000010101001101101101100 ; end 
      12'd85: begin cos_tmp = 24'b001111110001010011001101 ; sin_tmp = 24'b000010101100111000101011 ; end 
      12'd86: begin cos_tmp = 24'b001111110001010011001101 ; sin_tmp = 24'b000010101100111000101011 ; end 
      12'd87: begin cos_tmp = 24'b001111110000110000001000 ; sin_tmp = 24'b000010110000000011100011 ; end 
      12'd88: begin cos_tmp = 24'b001111110000001100011010 ; sin_tmp = 24'b000010110011001110010100 ; end 
      12'd89: begin cos_tmp = 24'b001111110000001100011010 ; sin_tmp = 24'b000010110011001110010100 ; end 
      12'd90: begin cos_tmp = 24'b001111101111101000000100 ; sin_tmp = 24'b000010110110011000111110 ; end 
      12'd91: begin cos_tmp = 24'b001111101111101000000100 ; sin_tmp = 24'b000010110110011000111110 ; end 
      12'd92: begin cos_tmp = 24'b001111101111000011000100 ; sin_tmp = 24'b000010111001100011100000 ; end 
      12'd93: begin cos_tmp = 24'b001111101110011101011100 ; sin_tmp = 24'b000010111100101101111011 ; end 
      12'd94: begin cos_tmp = 24'b001111101110011101011100 ; sin_tmp = 24'b000010111100101101111011 ; end 
      12'd95: begin cos_tmp = 24'b001111101101110111001011 ; sin_tmp = 24'b000010111111111000001110 ; end 
      12'd96: begin cos_tmp = 24'b001111101101110111001011 ; sin_tmp = 24'b000010111111111000001110 ; end 
      12'd97: begin cos_tmp = 24'b001111101101010000010010 ; sin_tmp = 24'b000011000011000010011010 ; end 
      12'd98: begin cos_tmp = 24'b001111101100101000110000 ; sin_tmp = 24'b000011000110001100011101 ; end 
      12'd99: begin cos_tmp = 24'b001111101100101000110000 ; sin_tmp = 24'b000011000110001100011101 ; end 
      12'd100: begin cos_tmp = 24'b001111101100000000100101 ; sin_tmp = 24'b000011001001010110011001 ; end 
      12'd101: begin cos_tmp = 24'b001111101011010111110010 ; sin_tmp = 24'b000011001100100000001100 ; end 
      12'd102: begin cos_tmp = 24'b001111101011010111110010 ; sin_tmp = 24'b000011001100100000001100 ; end 
      12'd103: begin cos_tmp = 24'b001111101010101110010110 ; sin_tmp = 24'b000011001111101001111000 ; end 
      12'd104: begin cos_tmp = 24'b001111101010101110010110 ; sin_tmp = 24'b000011001111101001111000 ; end 
      12'd105: begin cos_tmp = 24'b001111101010000100010010 ; sin_tmp = 24'b000011010010110011011010 ; end 
      12'd106: begin cos_tmp = 24'b001111101001011001100101 ; sin_tmp = 24'b000011010101111100110101 ; end 
      12'd107: begin cos_tmp = 24'b001111101001011001100101 ; sin_tmp = 24'b000011010101111100110101 ; end 
      12'd108: begin cos_tmp = 24'b001111101000101110010000 ; sin_tmp = 24'b000011011001000110000110 ; end 
      12'd109: begin cos_tmp = 24'b001111101000000010010010 ; sin_tmp = 24'b000011011100001111001111 ; end 
      12'd110: begin cos_tmp = 24'b001111101000000010010010 ; sin_tmp = 24'b000011011100001111001111 ; end 
      12'd111: begin cos_tmp = 24'b001111100111010101101100 ; sin_tmp = 24'b000011011111011000001111 ; end 
      12'd112: begin cos_tmp = 24'b001111100111010101101100 ; sin_tmp = 24'b000011011111011000001111 ; end 
      12'd113: begin cos_tmp = 24'b001111100110101000011101 ; sin_tmp = 24'b000011100010100001000110 ; end 
      12'd114: begin cos_tmp = 24'b001111100101111010100110 ; sin_tmp = 24'b000011100101101001110100 ; end 
      12'd115: begin cos_tmp = 24'b001111100101111010100110 ; sin_tmp = 24'b000011100101101001110100 ; end 
      12'd116: begin cos_tmp = 24'b001111100101001100000111 ; sin_tmp = 24'b000011101000110010011000 ; end 
      12'd117: begin cos_tmp = 24'b001111100100011100111111 ; sin_tmp = 24'b000011101011111010110011 ; end 
      12'd118: begin cos_tmp = 24'b001111100100011100111111 ; sin_tmp = 24'b000011101011111010110011 ; end 
      12'd119: begin cos_tmp = 24'b001111100011101101001111 ; sin_tmp = 24'b000011101111000011000101 ; end 
      12'd120: begin cos_tmp = 24'b001111100011101101001111 ; sin_tmp = 24'b000011101111000011000101 ; end 
      12'd121: begin cos_tmp = 24'b001111100010111100110111 ; sin_tmp = 24'b000011110010001011001101 ; end 
      12'd122: begin cos_tmp = 24'b001111100010001011110110 ; sin_tmp = 24'b000011110101010011001011 ; end 
      12'd123: begin cos_tmp = 24'b001111100010001011110110 ; sin_tmp = 24'b000011110101010011001011 ; end 
      12'd124: begin cos_tmp = 24'b001111100001011010001110 ; sin_tmp = 24'b000011111000011010111111 ; end 
      12'd125: begin cos_tmp = 24'b001111100000100111111101 ; sin_tmp = 24'b000011111011100010101001 ; end 
      12'd126: begin cos_tmp = 24'b001111100000100111111101 ; sin_tmp = 24'b000011111011100010101001 ; end 
      12'd127: begin cos_tmp = 24'b001111011111110101000100 ; sin_tmp = 24'b000011111110101010001001 ; end 
      12'd128: begin cos_tmp = 24'b001111011111110101000100 ; sin_tmp = 24'b000011111110101010001001 ; end 
      12'd129: begin cos_tmp = 24'b001111011111000001100011 ; sin_tmp = 24'b000100000001110001011111 ; end 
      12'd130: begin cos_tmp = 24'b001111011110001101011010 ; sin_tmp = 24'b000100000100111000101010 ; end 
      12'd131: begin cos_tmp = 24'b001111011110001101011010 ; sin_tmp = 24'b000100000100111000101010 ; end 
      12'd132: begin cos_tmp = 24'b001111011101011000101001 ; sin_tmp = 24'b000100000111111111101011 ; end 
      12'd133: begin cos_tmp = 24'b001111011101011000101001 ; sin_tmp = 24'b000100000111111111101011 ; end 
      12'd134: begin cos_tmp = 24'b001111011100100011010000 ; sin_tmp = 24'b000100001011000110100001 ; end 
      12'd135: begin cos_tmp = 24'b001111011011101101001111 ; sin_tmp = 24'b000100001110001101001100 ; end 
      12'd136: begin cos_tmp = 24'b001111011011101101001111 ; sin_tmp = 24'b000100001110001101001100 ; end 
      12'd137: begin cos_tmp = 24'b001111011010110110100110 ; sin_tmp = 24'b000100010001010011101100 ; end 
      12'd138: begin cos_tmp = 24'b001111011001111111010101 ; sin_tmp = 24'b000100010100011010000001 ; end 
      12'd139: begin cos_tmp = 24'b001111011001111111010101 ; sin_tmp = 24'b000100010100011010000001 ; end 
      12'd140: begin cos_tmp = 24'b001111011001000111011101 ; sin_tmp = 24'b000100010111100000001011 ; end 
      12'd141: begin cos_tmp = 24'b001111011001000111011101 ; sin_tmp = 24'b000100010111100000001011 ; end 
      12'd142: begin cos_tmp = 24'b001111011000001110111100 ; sin_tmp = 24'b000100011010100110001010 ; end 
      12'd143: begin cos_tmp = 24'b001111010111010101110100 ; sin_tmp = 24'b000100011101101011111110 ; end 
      12'd144: begin cos_tmp = 24'b001111010111010101110100 ; sin_tmp = 24'b000100011101101011111110 ; end 
      12'd145: begin cos_tmp = 24'b001111010110011100000100 ; sin_tmp = 24'b000100100000110001100101 ; end 
      12'd146: begin cos_tmp = 24'b001111010101100001101100 ; sin_tmp = 24'b000100100011110111000001 ; end 
      12'd147: begin cos_tmp = 24'b001111010101100001101100 ; sin_tmp = 24'b000100100011110111000001 ; end 
      12'd148: begin cos_tmp = 24'b001111010100100110101100 ; sin_tmp = 24'b000100100110111100010010 ; end 
      12'd149: begin cos_tmp = 24'b001111010100100110101100 ; sin_tmp = 24'b000100100110111100010010 ; end 
      12'd150: begin cos_tmp = 24'b001111010011101011000101 ; sin_tmp = 24'b000100101010000001010110 ; end 
      12'd151: begin cos_tmp = 24'b001111010010101110110110 ; sin_tmp = 24'b000100101101000110001111 ; end 
      12'd152: begin cos_tmp = 24'b001111010010101110110110 ; sin_tmp = 24'b000100101101000110001111 ; end 
      12'd153: begin cos_tmp = 24'b001111010001110010000000 ; sin_tmp = 24'b000100110000001010111011 ; end 
      12'd154: begin cos_tmp = 24'b001111010000110100100010 ; sin_tmp = 24'b000100110011001111011011 ; end 
      12'd155: begin cos_tmp = 24'b001111010000110100100010 ; sin_tmp = 24'b000100110011001111011011 ; end 
      12'd156: begin cos_tmp = 24'b001111001111110110011101 ; sin_tmp = 24'b000100110110010011101110 ; end 
      12'd157: begin cos_tmp = 24'b001111001111110110011101 ; sin_tmp = 24'b000100110110010011101110 ; end 
      12'd158: begin cos_tmp = 24'b001111001110110111110000 ; sin_tmp = 24'b000100111001010111110101 ; end 
      12'd159: begin cos_tmp = 24'b001111001101111000011100 ; sin_tmp = 24'b000100111100011011101111 ; end 
      12'd160: begin cos_tmp = 24'b001111001101111000011100 ; sin_tmp = 24'b000100111100011011101111 ; end 
      12'd161: begin cos_tmp = 24'b001111001100111000100001 ; sin_tmp = 24'b000100111111011111011101 ; end 
      12'd162: begin cos_tmp = 24'b001111001011110111111110 ; sin_tmp = 24'b000101000010100010111101 ; end 
      12'd163: begin cos_tmp = 24'b001111001011110111111110 ; sin_tmp = 24'b000101000010100010111101 ; end 
      12'd164: begin cos_tmp = 24'b001111001010110110110100 ; sin_tmp = 24'b000101000101100110010001 ; end 
      12'd165: begin cos_tmp = 24'b001111001010110110110100 ; sin_tmp = 24'b000101000101100110010001 ; end 
      12'd166: begin cos_tmp = 24'b001111001001110101000010 ; sin_tmp = 24'b000101001000101001010111 ; end 
      12'd167: begin cos_tmp = 24'b001111001000110010101010 ; sin_tmp = 24'b000101001011101100010000 ; end 
      12'd168: begin cos_tmp = 24'b001111001000110010101010 ; sin_tmp = 24'b000101001011101100010000 ; end 
      12'd169: begin cos_tmp = 24'b001111000111101111101010 ; sin_tmp = 24'b000101001110101110111100 ; end 
      12'd170: begin cos_tmp = 24'b001111000111101111101010 ; sin_tmp = 24'b000101001110101110111100 ; end 
      12'd171: begin cos_tmp = 24'b001111000110101100000011 ; sin_tmp = 24'b000101010001110001011010 ; end 
      12'd172: begin cos_tmp = 24'b001111000101100111110101 ; sin_tmp = 24'b000101010100110011101010 ; end 
      12'd173: begin cos_tmp = 24'b001111000101100111110101 ; sin_tmp = 24'b000101010100110011101010 ; end 
      12'd174: begin cos_tmp = 24'b001111000100100011000000 ; sin_tmp = 24'b000101010111110101101101 ; end 
      12'd175: begin cos_tmp = 24'b001111000011011101100100 ; sin_tmp = 24'b000101011010110111100010 ; end 
      12'd176: begin cos_tmp = 24'b001111000011011101100100 ; sin_tmp = 24'b000101011010110111100010 ; end 
      12'd177: begin cos_tmp = 24'b001111000010010111100001 ; sin_tmp = 24'b000101011101111001001001 ; end 
      12'd178: begin cos_tmp = 24'b001111000010010111100001 ; sin_tmp = 24'b000101011101111001001001 ; end 
      12'd179: begin cos_tmp = 24'b001111000001010000110111 ; sin_tmp = 24'b000101100000111010100001 ; end 
      12'd180: begin cos_tmp = 24'b001111000000001001100110 ; sin_tmp = 24'b000101100011111011101100 ; end 
      12'd181: begin cos_tmp = 24'b001111000000001001100110 ; sin_tmp = 24'b000101100011111011101100 ; end 
      12'd182: begin cos_tmp = 24'b001110111111000001101111 ; sin_tmp = 24'b000101100110111100101000 ; end 
      12'd183: begin cos_tmp = 24'b001110111101111001010001 ; sin_tmp = 24'b000101101001111101010101 ; end 
      12'd184: begin cos_tmp = 24'b001110111101111001010001 ; sin_tmp = 24'b000101101001111101010101 ; end 
      12'd185: begin cos_tmp = 24'b001110111100110000001100 ; sin_tmp = 24'b000101101100111101110100 ; end 
      12'd186: begin cos_tmp = 24'b001110111100110000001100 ; sin_tmp = 24'b000101101100111101110100 ; end 
      12'd187: begin cos_tmp = 24'b001110111011100110100000 ; sin_tmp = 24'b000101101111111110000100 ; end 
      12'd188: begin cos_tmp = 24'b001110111010011100001110 ; sin_tmp = 24'b000101110010111110000101 ; end 
      12'd189: begin cos_tmp = 24'b001110111010011100001110 ; sin_tmp = 24'b000101110010111110000101 ; end 
      12'd190: begin cos_tmp = 24'b001110111001010001010101 ; sin_tmp = 24'b000101110101111101110111 ; end 
      12'd191: begin cos_tmp = 24'b001110111000000101110101 ; sin_tmp = 24'b000101111000111101011010 ; end 
      12'd192: begin cos_tmp = 24'b001110111000000101110101 ; sin_tmp = 24'b000101111000111101011010 ; end 
      12'd193: begin cos_tmp = 24'b001110110110111001101111 ; sin_tmp = 24'b000101111011111100101110 ; end 
      12'd194: begin cos_tmp = 24'b001110110110111001101111 ; sin_tmp = 24'b000101111011111100101110 ; end 
      12'd195: begin cos_tmp = 24'b001110110101101101000011 ; sin_tmp = 24'b000101111110111011110011 ; end 
      12'd196: begin cos_tmp = 24'b001110110100011111110000 ; sin_tmp = 24'b000110000001111010101000 ; end 
      12'd197: begin cos_tmp = 24'b001110110100011111110000 ; sin_tmp = 24'b000110000001111010101000 ; end 
      12'd198: begin cos_tmp = 24'b001110110011010001110111 ; sin_tmp = 24'b000110000100111001001101 ; end 
      12'd199: begin cos_tmp = 24'b001110110010000011011000 ; sin_tmp = 24'b000110000111110111100011 ; end 
      12'd200: begin cos_tmp = 24'b001110110010000011011000 ; sin_tmp = 24'b000110000111110111100011 ; end 
      12'd201: begin cos_tmp = 24'b001110110000110100010010 ; sin_tmp = 24'b000110001010110101101000 ; end 
      12'd202: begin cos_tmp = 24'b001110110000110100010010 ; sin_tmp = 24'b000110001010110101101000 ; end 
      12'd203: begin cos_tmp = 24'b001110101111100100100110 ; sin_tmp = 24'b000110001101110011011110 ; end 
      12'd204: begin cos_tmp = 24'b001110101110010100010100 ; sin_tmp = 24'b000110010000110001000100 ; end 
      12'd205: begin cos_tmp = 24'b001110101110010100010100 ; sin_tmp = 24'b000110010000110001000100 ; end 
      12'd206: begin cos_tmp = 24'b001110101101000011011100 ; sin_tmp = 24'b000110010011101110011010 ; end 
      12'd207: begin cos_tmp = 24'b001110101011110001111110 ; sin_tmp = 24'b000110010110101011011111 ; end 
      12'd208: begin cos_tmp = 24'b001110101011110001111110 ; sin_tmp = 24'b000110010110101011011111 ; end 
      12'd209: begin cos_tmp = 24'b001110101010011111111010 ; sin_tmp = 24'b000110011001101000010100 ; end 
      12'd210: begin cos_tmp = 24'b001110101010011111111010 ; sin_tmp = 24'b000110011001101000010100 ; end 
      12'd211: begin cos_tmp = 24'b001110101001001101010000 ; sin_tmp = 24'b000110011100100100111000 ; end 
      12'd212: begin cos_tmp = 24'b001110100111111010000000 ; sin_tmp = 24'b000110011111100001001100 ; end 
      12'd213: begin cos_tmp = 24'b001110100111111010000000 ; sin_tmp = 24'b000110011111100001001100 ; end 
      12'd214: begin cos_tmp = 24'b001110100110100110001010 ; sin_tmp = 24'b000110100010011101001110 ; end 
      12'd215: begin cos_tmp = 24'b001110100110100110001010 ; sin_tmp = 24'b000110100010011101001110 ; end 
      12'd216: begin cos_tmp = 24'b001110100101010001101110 ; sin_tmp = 24'b000110100101011001000000 ; end 
      12'd217: begin cos_tmp = 24'b001110100011111100101101 ; sin_tmp = 24'b000110101000010100100001 ; end 
      12'd218: begin cos_tmp = 24'b001110100011111100101101 ; sin_tmp = 24'b000110101000010100100001 ; end 
      12'd219: begin cos_tmp = 24'b001110100010100111000110 ; sin_tmp = 24'b000110101011001111110001 ; end 
      12'd220: begin cos_tmp = 24'b001110100001010000111010 ; sin_tmp = 24'b000110101110001010101111 ; end 
      12'd221: begin cos_tmp = 24'b001110100001010000111010 ; sin_tmp = 24'b000110101110001010101111 ; end 
      12'd222: begin cos_tmp = 24'b001110011111111010000111 ; sin_tmp = 24'b000110110001000101011100 ; end 
      12'd223: begin cos_tmp = 24'b001110011111111010000111 ; sin_tmp = 24'b000110110001000101011100 ; end 
      12'd224: begin cos_tmp = 24'b001110011110100010110000 ; sin_tmp = 24'b000110110011111111111000 ; end 
      12'd225: begin cos_tmp = 24'b001110011101001010110011 ; sin_tmp = 24'b000110110110111010000010 ; end 
      12'd226: begin cos_tmp = 24'b001110011101001010110011 ; sin_tmp = 24'b000110110110111010000010 ; end 
      12'd227: begin cos_tmp = 24'b001110011011110010010000 ; sin_tmp = 24'b000110111001110011111010 ; end 
      12'd228: begin cos_tmp = 24'b001110011010011001001000 ; sin_tmp = 24'b000110111100101101100000 ; end 
      12'd229: begin cos_tmp = 24'b001110011010011001001000 ; sin_tmp = 24'b000110111100101101100000 ; end 
      12'd230: begin cos_tmp = 24'b001110011000111111011011 ; sin_tmp = 24'b000110111111100110110100 ; end 
      12'd231: begin cos_tmp = 24'b001110011000111111011011 ; sin_tmp = 24'b000110111111100110110100 ; end 
      12'd232: begin cos_tmp = 24'b001110010111100101001001 ; sin_tmp = 24'b000111000010011111110111 ; end 
      12'd233: begin cos_tmp = 24'b001110010110001010010001 ; sin_tmp = 24'b000111000101011000100111 ; end 
      12'd234: begin cos_tmp = 24'b001110010110001010010001 ; sin_tmp = 24'b000111000101011000100111 ; end 
      12'd235: begin cos_tmp = 24'b001110010100101110110100 ; sin_tmp = 24'b000111001000010001000100 ; end 
      12'd236: begin cos_tmp = 24'b001110010011010010110011 ; sin_tmp = 24'b000111001011001001010000 ; end 
      12'd237: begin cos_tmp = 24'b001110010011010010110011 ; sin_tmp = 24'b000111001011001001010000 ; end 
      12'd238: begin cos_tmp = 24'b001110010001110110001100 ; sin_tmp = 24'b000111001110000001001000 ; end 
      12'd239: begin cos_tmp = 24'b001110010001110110001100 ; sin_tmp = 24'b000111001110000001001000 ; end 
      12'd240: begin cos_tmp = 24'b001110010000011001000000 ; sin_tmp = 24'b000111010000111000101110 ; end 
      12'd241: begin cos_tmp = 24'b001110001110111011010000 ; sin_tmp = 24'b000111010011110000000001 ; end 
      12'd242: begin cos_tmp = 24'b001110001110111011010000 ; sin_tmp = 24'b000111010011110000000001 ; end 
      12'd243: begin cos_tmp = 24'b001110001101011100111010 ; sin_tmp = 24'b000111010110100111000010 ; end 
      12'd244: begin cos_tmp = 24'b001110001011111110000000 ; sin_tmp = 24'b000111011001011101101111 ; end 
      12'd245: begin cos_tmp = 24'b001110001011111110000000 ; sin_tmp = 24'b000111011001011101101111 ; end 
      12'd246: begin cos_tmp = 24'b001110001010011110100001 ; sin_tmp = 24'b000111011100010100001001 ; end 
      12'd247: begin cos_tmp = 24'b001110001010011110100001 ; sin_tmp = 24'b000111011100010100001001 ; end 
      12'd248: begin cos_tmp = 24'b001110001000111110011110 ; sin_tmp = 24'b000111011111001010010000 ; end 
      12'd249: begin cos_tmp = 24'b001110000111011101110110 ; sin_tmp = 24'b000111100010000000000011 ; end 
      12'd250: begin cos_tmp = 24'b001110000111011101110110 ; sin_tmp = 24'b000111100010000000000011 ; end 
      12'd251: begin cos_tmp = 24'b001110000101111100101001 ; sin_tmp = 24'b000111100100110101100011 ; end 
      12'd252: begin cos_tmp = 24'b001110000101111100101001 ; sin_tmp = 24'b000111100100110101100011 ; end 
      12'd253: begin cos_tmp = 24'b001110000100011010111000 ; sin_tmp = 24'b000111100111101010110000 ; end 
      12'd254: begin cos_tmp = 24'b001110000010111000100010 ; sin_tmp = 24'b000111101010011111101000 ; end 
      12'd255: begin cos_tmp = 24'b001110000010111000100010 ; sin_tmp = 24'b000111101010011111101000 ; end 
      12'd256: begin cos_tmp = 24'b001110000001010101101001 ; sin_tmp = 24'b000111101101010100001101 ; end 
      12'd257: begin cos_tmp = 24'b001101111111110010001011 ; sin_tmp = 24'b000111110000001000011110 ; end 
      12'd258: begin cos_tmp = 24'b001101111111110010001011 ; sin_tmp = 24'b000111110000001000011110 ; end 
      12'd259: begin cos_tmp = 24'b001101111110001110001000 ; sin_tmp = 24'b000111110010111100011011 ; end 
      12'd260: begin cos_tmp = 24'b001101111110001110001000 ; sin_tmp = 24'b000111110010111100011011 ; end 
      12'd261: begin cos_tmp = 24'b001101111100101001100010 ; sin_tmp = 24'b000111110101110000000100 ; end 
      12'd262: begin cos_tmp = 24'b001101111011000100010111 ; sin_tmp = 24'b000111111000100011011000 ; end 
      12'd263: begin cos_tmp = 24'b001101111011000100010111 ; sin_tmp = 24'b000111111000100011011000 ; end 
      12'd264: begin cos_tmp = 24'b001101111001011110101001 ; sin_tmp = 24'b000111111011010110011000 ; end 
      12'd265: begin cos_tmp = 24'b001101110111111000010110 ; sin_tmp = 24'b000111111110001001000100 ; end 
      12'd266: begin cos_tmp = 24'b001101110111111000010110 ; sin_tmp = 24'b000111111110001001000100 ; end 
      12'd267: begin cos_tmp = 24'b001101110110010001100000 ; sin_tmp = 24'b001000000000111011011011 ; end 
      12'd268: begin cos_tmp = 24'b001101110110010001100000 ; sin_tmp = 24'b001000000000111011011011 ; end 
      12'd269: begin cos_tmp = 24'b001101110100101010000101 ; sin_tmp = 24'b001000000011101101011101 ; end 
      12'd270: begin cos_tmp = 24'b001101110011000010000111 ; sin_tmp = 24'b001000000110011111001010 ; end 
      12'd271: begin cos_tmp = 24'b001101110011000010000111 ; sin_tmp = 24'b001000000110011111001010 ; end 
      12'd272: begin cos_tmp = 24'b001101110001011001100110 ; sin_tmp = 24'b001000001001010000100010 ; end 
      12'd273: begin cos_tmp = 24'b001101101111110000100000 ; sin_tmp = 24'b001000001100000001100110 ; end 
      12'd274: begin cos_tmp = 24'b001101101111110000100000 ; sin_tmp = 24'b001000001100000001100110 ; end 
      12'd275: begin cos_tmp = 24'b001101101110000110110111 ; sin_tmp = 24'b001000001110110010010100 ; end 
      12'd276: begin cos_tmp = 24'b001101101110000110110111 ; sin_tmp = 24'b001000001110110010010100 ; end 
      12'd277: begin cos_tmp = 24'b001101101100011100101011 ; sin_tmp = 24'b001000010001100010101101 ; end 
      12'd278: begin cos_tmp = 24'b001101101010110001111011 ; sin_tmp = 24'b001000010100010010110000 ; end 
      12'd279: begin cos_tmp = 24'b001101101010110001111011 ; sin_tmp = 24'b001000010100010010110000 ; end 
      12'd280: begin cos_tmp = 24'b001101101001000110101000 ; sin_tmp = 24'b001000010111000010011110 ; end 
      12'd281: begin cos_tmp = 24'b001101100111011010110010 ; sin_tmp = 24'b001000011001110001110110 ; end 
      12'd282: begin cos_tmp = 24'b001101100111011010110010 ; sin_tmp = 24'b001000011001110001110110 ; end 
      12'd283: begin cos_tmp = 24'b001101100101101110011000 ; sin_tmp = 24'b001000011100100000111001 ; end 
      12'd284: begin cos_tmp = 24'b001101100101101110011000 ; sin_tmp = 24'b001000011100100000111001 ; end 
      12'd285: begin cos_tmp = 24'b001101100100000001011011 ; sin_tmp = 24'b001000011111001111100101 ; end 
      12'd286: begin cos_tmp = 24'b001101100010010011111011 ; sin_tmp = 24'b001000100001111101111100 ; end 
      12'd287: begin cos_tmp = 24'b001101100010010011111011 ; sin_tmp = 24'b001000100001111101111100 ; end 
      12'd288: begin cos_tmp = 24'b001101100000100101111000 ; sin_tmp = 24'b001000100100101011111100 ; end 
      12'd289: begin cos_tmp = 24'b001101100000100101111000 ; sin_tmp = 24'b001000100100101011111100 ; end 
      12'd290: begin cos_tmp = 24'b001101011110110111010010 ; sin_tmp = 24'b001000100111011001100111 ; end 
      12'd291: begin cos_tmp = 24'b001101011101001000001001 ; sin_tmp = 24'b001000101010000110111011 ; end 
      12'd292: begin cos_tmp = 24'b001101011101001000001001 ; sin_tmp = 24'b001000101010000110111011 ; end 
      12'd293: begin cos_tmp = 24'b001101011011011000011110 ; sin_tmp = 24'b001000101100110011111001 ; end 
      12'd294: begin cos_tmp = 24'b001101011001101000001111 ; sin_tmp = 24'b001000101111100000100000 ; end 
      12'd295: begin cos_tmp = 24'b001101011001101000001111 ; sin_tmp = 24'b001000101111100000100000 ; end 
      12'd296: begin cos_tmp = 24'b001101010111110111011110 ; sin_tmp = 24'b001000110010001100110001 ; end 
      12'd297: begin cos_tmp = 24'b001101010111110111011110 ; sin_tmp = 24'b001000110010001100110001 ; end 
      12'd298: begin cos_tmp = 24'b001101010110000110001011 ; sin_tmp = 24'b001000110100111000101010 ; end 
      12'd299: begin cos_tmp = 24'b001101010100010100010100 ; sin_tmp = 24'b001000110111100100001110 ; end 
      12'd300: begin cos_tmp = 24'b001101010100010100010100 ; sin_tmp = 24'b001000110111100100001110 ; end 
      12'd301: begin cos_tmp = 24'b001101010010100001111100 ; sin_tmp = 24'b001000111010001111011010 ; end 
      12'd302: begin cos_tmp = 24'b001101010000101111000001 ; sin_tmp = 24'b001000111100111010001111 ; end 
      12'd303: begin cos_tmp = 24'b001101010000101111000001 ; sin_tmp = 24'b001000111100111010001111 ; end 
      12'd304: begin cos_tmp = 24'b001101001110111011100011 ; sin_tmp = 24'b001000111111100100101101 ; end 
      12'd305: begin cos_tmp = 24'b001101001110111011100011 ; sin_tmp = 24'b001000111111100100101101 ; end 
      12'd306: begin cos_tmp = 24'b001101001101000111100100 ; sin_tmp = 24'b001001000010001110110011 ; end 
      12'd307: begin cos_tmp = 24'b001101001011010011000010 ; sin_tmp = 24'b001001000100111000100010 ; end 
      12'd308: begin cos_tmp = 24'b001101001011010011000010 ; sin_tmp = 24'b001001000100111000100010 ; end 
      12'd309: begin cos_tmp = 24'b001101001001011101111110 ; sin_tmp = 24'b001001000111100001111010 ; end 
      12'd310: begin cos_tmp = 24'b001101000111101000011000 ; sin_tmp = 24'b001001001010001010111010 ; end 
      12'd311: begin cos_tmp = 24'b001101000111101000011000 ; sin_tmp = 24'b001001001010001010111010 ; end 
      12'd312: begin cos_tmp = 24'b001101000101110010010001 ; sin_tmp = 24'b001001001100110011100011 ; end 
      12'd313: begin cos_tmp = 24'b001101000101110010010001 ; sin_tmp = 24'b001001001100110011100011 ; end 
      12'd314: begin cos_tmp = 24'b001101000011111011100111 ; sin_tmp = 24'b001001001111011011110100 ; end 
      12'd315: begin cos_tmp = 24'b001101000010000100011100 ; sin_tmp = 24'b001001010010000011101100 ; end 
      12'd316: begin cos_tmp = 24'b001101000010000100011100 ; sin_tmp = 24'b001001010010000011101100 ; end 
      12'd317: begin cos_tmp = 24'b001101000000001100101110 ; sin_tmp = 24'b001001010100101011001101 ; end 
      12'd318: begin cos_tmp = 24'b001100111110010100100000 ; sin_tmp = 24'b001001010111010010010110 ; end 
      12'd319: begin cos_tmp = 24'b001100111110010100100000 ; sin_tmp = 24'b001001010111010010010110 ; end 
      12'd320: begin cos_tmp = 24'b001100111100011011101111 ; sin_tmp = 24'b001001011001111001000110 ; end 
      12'd321: begin cos_tmp = 24'b001100111100011011101111 ; sin_tmp = 24'b001001011001111001000110 ; end 
      12'd322: begin cos_tmp = 24'b001100111010100010011101 ; sin_tmp = 24'b001001011100011111011110 ; end 
      12'd323: begin cos_tmp = 24'b001100111000101000101010 ; sin_tmp = 24'b001001011111000101011110 ; end 
      12'd324: begin cos_tmp = 24'b001100111000101000101010 ; sin_tmp = 24'b001001011111000101011110 ; end 
      12'd325: begin cos_tmp = 24'b001100110110101110010101 ; sin_tmp = 24'b001001100001101011000101 ; end 
      12'd326: begin cos_tmp = 24'b001100110110101110010101 ; sin_tmp = 24'b001001100001101011000101 ; end 
      12'd327: begin cos_tmp = 24'b001100110100110011100000 ; sin_tmp = 24'b001001100100010000010011 ; end 
      12'd328: begin cos_tmp = 24'b001100110010111000001001 ; sin_tmp = 24'b001001100110110101001001 ; end 
      12'd329: begin cos_tmp = 24'b001100110010111000001001 ; sin_tmp = 24'b001001100110110101001001 ; end 
      12'd330: begin cos_tmp = 24'b001100110000111100010000 ; sin_tmp = 24'b001001101001011001100110 ; end 
      12'd331: begin cos_tmp = 24'b001100101110111111110111 ; sin_tmp = 24'b001001101011111101101010 ; end 
      12'd332: begin cos_tmp = 24'b001100101110111111110111 ; sin_tmp = 24'b001001101011111101101010 ; end 
      12'd333: begin cos_tmp = 24'b001100101101000010111101 ; sin_tmp = 24'b001001101110100001010100 ; end 
      12'd334: begin cos_tmp = 24'b001100101101000010111101 ; sin_tmp = 24'b001001101110100001010100 ; end 
      12'd335: begin cos_tmp = 24'b001100101011000101100010 ; sin_tmp = 24'b001001110001000100100110 ; end 
      12'd336: begin cos_tmp = 24'b001100101001000111100110 ; sin_tmp = 24'b001001110011100111011111 ; end 
      12'd337: begin cos_tmp = 24'b001100101001000111100110 ; sin_tmp = 24'b001001110011100111011111 ; end 
      12'd338: begin cos_tmp = 24'b001100100111001001001010 ; sin_tmp = 24'b001001110110001001111110 ; end 
      12'd339: begin cos_tmp = 24'b001100100101001010001101 ; sin_tmp = 24'b001001111000101100000011 ; end 
      12'd340: begin cos_tmp = 24'b001100100101001010001101 ; sin_tmp = 24'b001001111000101100000011 ; end 
      12'd341: begin cos_tmp = 24'b001100100011001010101111 ; sin_tmp = 24'b001001111011001101101111 ; end 
      12'd342: begin cos_tmp = 24'b001100100011001010101111 ; sin_tmp = 24'b001001111011001101101111 ; end 
      12'd343: begin cos_tmp = 24'b001100100001001010110001 ; sin_tmp = 24'b001001111101101111000001 ; end 
      12'd344: begin cos_tmp = 24'b001100011111001010010010 ; sin_tmp = 24'b001010000000001111111010 ; end 
      12'd345: begin cos_tmp = 24'b001100011111001010010010 ; sin_tmp = 24'b001010000000001111111010 ; end 
      12'd346: begin cos_tmp = 24'b001100011101001001010100 ; sin_tmp = 24'b001010000010110000011000 ; end 
      12'd347: begin cos_tmp = 24'b001100011011000111110100 ; sin_tmp = 24'b001010000101010000011101 ; end 
      12'd348: begin cos_tmp = 24'b001100011011000111110100 ; sin_tmp = 24'b001010000101010000011101 ; end 
      12'd349: begin cos_tmp = 24'b001100011001000101110101 ; sin_tmp = 24'b001010000111110000001000 ; end 
      12'd350: begin cos_tmp = 24'b001100011001000101110101 ; sin_tmp = 24'b001010000111110000001000 ; end 
      12'd351: begin cos_tmp = 24'b001100010111000011010110 ; sin_tmp = 24'b001010001010001111011000 ; end 
      12'd352: begin cos_tmp = 24'b001100010101000000010111 ; sin_tmp = 24'b001010001100101110001110 ; end 
      12'd353: begin cos_tmp = 24'b001100010101000000010111 ; sin_tmp = 24'b001010001100101110001110 ; end 
      12'd354: begin cos_tmp = 24'b001100010010111100111000 ; sin_tmp = 24'b001010001111001100101010 ; end 
      12'd355: begin cos_tmp = 24'b001100010000111000111001 ; sin_tmp = 24'b001010010001101010101011 ; end 
      12'd356: begin cos_tmp = 24'b001100010000111000111001 ; sin_tmp = 24'b001010010001101010101011 ; end 
      12'd357: begin cos_tmp = 24'b001100001110110100011010 ; sin_tmp = 24'b001010010100001000010001 ; end 
      12'd358: begin cos_tmp = 24'b001100001110110100011010 ; sin_tmp = 24'b001010010100001000010001 ; end 
      12'd359: begin cos_tmp = 24'b001100001100101111011100 ; sin_tmp = 24'b001010010110100101011101 ; end 
      12'd360: begin cos_tmp = 24'b001100001010101001111110 ; sin_tmp = 24'b001010011001000010001111 ; end 
      12'd361: begin cos_tmp = 24'b001100001010101001111110 ; sin_tmp = 24'b001010011001000010001111 ; end 
      12'd362: begin cos_tmp = 24'b001100001000100100000000 ; sin_tmp = 24'b001010011011011110100101 ; end 
      12'd363: begin cos_tmp = 24'b001100001000100100000000 ; sin_tmp = 24'b001010011011011110100101 ; end 
      12'd364: begin cos_tmp = 24'b001100000110011101100100 ; sin_tmp = 24'b001010011101111010100000 ; end 
      12'd365: begin cos_tmp = 24'b001100000100010110101000 ; sin_tmp = 24'b001010100000010110000000 ; end 
      12'd366: begin cos_tmp = 24'b001100000100010110101000 ; sin_tmp = 24'b001010100000010110000000 ; end 
      12'd367: begin cos_tmp = 24'b001100000010001111001100 ; sin_tmp = 24'b001010100010110001000101 ; end 
      12'd368: begin cos_tmp = 24'b001100000000000111010010 ; sin_tmp = 24'b001010100101001011101111 ; end 
      12'd369: begin cos_tmp = 24'b001100000000000111010010 ; sin_tmp = 24'b001010100101001011101111 ; end 
      12'd370: begin cos_tmp = 24'b001011111101111110111000 ; sin_tmp = 24'b001010100111100101111101 ; end 
      12'd371: begin cos_tmp = 24'b001011111101111110111000 ; sin_tmp = 24'b001010100111100101111101 ; end 
      12'd372: begin cos_tmp = 24'b001011111011110110000000 ; sin_tmp = 24'b001010101001111111110000 ; end 
      12'd373: begin cos_tmp = 24'b001011111001101100101001 ; sin_tmp = 24'b001010101100011001001000 ; end 
      12'd374: begin cos_tmp = 24'b001011111001101100101001 ; sin_tmp = 24'b001010101100011001001000 ; end 
      12'd375: begin cos_tmp = 24'b001011110111100010110010 ; sin_tmp = 24'b001010101110110010000011 ; end 
      12'd376: begin cos_tmp = 24'b001011110101011000011110 ; sin_tmp = 24'b001010110001001010100011 ; end 
      12'd377: begin cos_tmp = 24'b001011110101011000011110 ; sin_tmp = 24'b001010110001001010100011 ; end 
      12'd378: begin cos_tmp = 24'b001011110011001101101010 ; sin_tmp = 24'b001010110011100010100111 ; end 
      12'd379: begin cos_tmp = 24'b001011110011001101101010 ; sin_tmp = 24'b001010110011100010100111 ; end 
      12'd380: begin cos_tmp = 24'b001011110001000010011000 ; sin_tmp = 24'b001010110101111010001111 ; end 
      12'd381: begin cos_tmp = 24'b001011101110110110101000 ; sin_tmp = 24'b001010111000010001011011 ; end 
      12'd382: begin cos_tmp = 24'b001011101110110110101000 ; sin_tmp = 24'b001010111000010001011011 ; end 
      12'd383: begin cos_tmp = 24'b001011101100101010011001 ; sin_tmp = 24'b001010111010101000001011 ; end 
      12'd384: begin cos_tmp = 24'b001011101010011101101100 ; sin_tmp = 24'b001010111100111110011111 ; end 
      12'd385: begin cos_tmp = 24'b001011101010011101101100 ; sin_tmp = 24'b001010111100111110011111 ; end 
      12'd386: begin cos_tmp = 24'b001011101000010000100001 ; sin_tmp = 24'b001010111111010100010110 ; end 
      12'd387: begin cos_tmp = 24'b001011101000010000100001 ; sin_tmp = 24'b001010111111010100010110 ; end 
      12'd388: begin cos_tmp = 24'b001011100110000010111000 ; sin_tmp = 24'b001011000001101001110001 ; end 
      12'd389: begin cos_tmp = 24'b001011100011110100110000 ; sin_tmp = 24'b001011000011111110101111 ; end 
      12'd390: begin cos_tmp = 24'b001011100011110100110000 ; sin_tmp = 24'b001011000011111110101111 ; end 
      12'd391: begin cos_tmp = 24'b001011100001100110001011 ; sin_tmp = 24'b001011000110010011010001 ; end 
      12'd392: begin cos_tmp = 24'b001011011111010111001000 ; sin_tmp = 24'b001011001000100111010110 ; end 
      12'd393: begin cos_tmp = 24'b001011011111010111001000 ; sin_tmp = 24'b001011001000100111010110 ; end 
      12'd394: begin cos_tmp = 24'b001011011101000111100111 ; sin_tmp = 24'b001011001010111010111110 ; end 
      12'd395: begin cos_tmp = 24'b001011011101000111100111 ; sin_tmp = 24'b001011001010111010111110 ; end 
      12'd396: begin cos_tmp = 24'b001011011010110111101001 ; sin_tmp = 24'b001011001101001110001001 ; end 
      12'd397: begin cos_tmp = 24'b001011011000100111001101 ; sin_tmp = 24'b001011001111100000111000 ; end 
      12'd398: begin cos_tmp = 24'b001011011000100111001101 ; sin_tmp = 24'b001011001111100000111000 ; end 
      12'd399: begin cos_tmp = 24'b001011010110010110010100 ; sin_tmp = 24'b001011010001110011001001 ; end 
      12'd400: begin cos_tmp = 24'b001011010110010110010100 ; sin_tmp = 24'b001011010001110011001001 ; end 
      12'd401: begin cos_tmp = 24'b001011010100000100111101 ; sin_tmp = 24'b001011010100000100111101 ; end 
      12'd402: begin cos_tmp = 24'b001011010001110011001001 ; sin_tmp = 24'b001011010110010110010100 ; end 
      12'd403: begin cos_tmp = 24'b001011010001110011001001 ; sin_tmp = 24'b001011010110010110010100 ; end 
      12'd404: begin cos_tmp = 24'b001011001111100000111000 ; sin_tmp = 24'b001011011000100111001101 ; end 
      12'd405: begin cos_tmp = 24'b001011001101001110001001 ; sin_tmp = 24'b001011011010110111101001 ; end 
      12'd406: begin cos_tmp = 24'b001011001101001110001001 ; sin_tmp = 24'b001011011010110111101001 ; end 
      12'd407: begin cos_tmp = 24'b001011001010111010111110 ; sin_tmp = 24'b001011011101000111100111 ; end 
      12'd408: begin cos_tmp = 24'b001011001010111010111110 ; sin_tmp = 24'b001011011101000111100111 ; end 
      12'd409: begin cos_tmp = 24'b001011001000100111010110 ; sin_tmp = 24'b001011011111010111001000 ; end 
      12'd410: begin cos_tmp = 24'b001011000110010011010001 ; sin_tmp = 24'b001011100001100110001011 ; end 
      12'd411: begin cos_tmp = 24'b001011000110010011010001 ; sin_tmp = 24'b001011100001100110001011 ; end 
      12'd412: begin cos_tmp = 24'b001011000011111110101111 ; sin_tmp = 24'b001011100011110100110000 ; end 
      12'd413: begin cos_tmp = 24'b001011000001101001110001 ; sin_tmp = 24'b001011100110000010111000 ; end 
      12'd414: begin cos_tmp = 24'b001011000001101001110001 ; sin_tmp = 24'b001011100110000010111000 ; end 
      12'd415: begin cos_tmp = 24'b001010111111010100010110 ; sin_tmp = 24'b001011101000010000100001 ; end 
      12'd416: begin cos_tmp = 24'b001010111111010100010110 ; sin_tmp = 24'b001011101000010000100001 ; end 
      12'd417: begin cos_tmp = 24'b001010111100111110011111 ; sin_tmp = 24'b001011101010011101101100 ; end 
      12'd418: begin cos_tmp = 24'b001010111010101000001011 ; sin_tmp = 24'b001011101100101010011001 ; end 
      12'd419: begin cos_tmp = 24'b001010111010101000001011 ; sin_tmp = 24'b001011101100101010011001 ; end 
      12'd420: begin cos_tmp = 24'b001010111000010001011011 ; sin_tmp = 24'b001011101110110110101000 ; end 
      12'd421: begin cos_tmp = 24'b001010110101111010001111 ; sin_tmp = 24'b001011110001000010011000 ; end 
      12'd422: begin cos_tmp = 24'b001010110101111010001111 ; sin_tmp = 24'b001011110001000010011000 ; end 
      12'd423: begin cos_tmp = 24'b001010110011100010100111 ; sin_tmp = 24'b001011110011001101101010 ; end 
      12'd424: begin cos_tmp = 24'b001010110011100010100111 ; sin_tmp = 24'b001011110011001101101010 ; end 
      12'd425: begin cos_tmp = 24'b001010110001001010100011 ; sin_tmp = 24'b001011110101011000011110 ; end 
      12'd426: begin cos_tmp = 24'b001010101110110010000011 ; sin_tmp = 24'b001011110111100010110010 ; end 
      12'd427: begin cos_tmp = 24'b001010101110110010000011 ; sin_tmp = 24'b001011110111100010110010 ; end 
      12'd428: begin cos_tmp = 24'b001010101100011001001000 ; sin_tmp = 24'b001011111001101100101001 ; end 
      12'd429: begin cos_tmp = 24'b001010101001111111110000 ; sin_tmp = 24'b001011111011110110000000 ; end 
      12'd430: begin cos_tmp = 24'b001010101001111111110000 ; sin_tmp = 24'b001011111011110110000000 ; end 
      12'd431: begin cos_tmp = 24'b001010100111100101111101 ; sin_tmp = 24'b001011111101111110111000 ; end 
      12'd432: begin cos_tmp = 24'b001010100111100101111101 ; sin_tmp = 24'b001011111101111110111000 ; end 
      12'd433: begin cos_tmp = 24'b001010100101001011101111 ; sin_tmp = 24'b001100000000000111010010 ; end 
      12'd434: begin cos_tmp = 24'b001010100010110001000101 ; sin_tmp = 24'b001100000010001111001100 ; end 
      12'd435: begin cos_tmp = 24'b001010100010110001000101 ; sin_tmp = 24'b001100000010001111001100 ; end 
      12'd436: begin cos_tmp = 24'b001010100000010110000000 ; sin_tmp = 24'b001100000100010110101000 ; end 
      12'd437: begin cos_tmp = 24'b001010100000010110000000 ; sin_tmp = 24'b001100000100010110101000 ; end 
      12'd438: begin cos_tmp = 24'b001010011101111010100000 ; sin_tmp = 24'b001100000110011101100100 ; end 
      12'd439: begin cos_tmp = 24'b001010011011011110100101 ; sin_tmp = 24'b001100001000100100000000 ; end 
      12'd440: begin cos_tmp = 24'b001010011011011110100101 ; sin_tmp = 24'b001100001000100100000000 ; end 
      12'd441: begin cos_tmp = 24'b001010011001000010001111 ; sin_tmp = 24'b001100001010101001111110 ; end 
      12'd442: begin cos_tmp = 24'b001010010110100101011101 ; sin_tmp = 24'b001100001100101111011100 ; end 
      12'd443: begin cos_tmp = 24'b001010010110100101011101 ; sin_tmp = 24'b001100001100101111011100 ; end 
      12'd444: begin cos_tmp = 24'b001010010100001000010001 ; sin_tmp = 24'b001100001110110100011010 ; end 
      12'd445: begin cos_tmp = 24'b001010010100001000010001 ; sin_tmp = 24'b001100001110110100011010 ; end 
      12'd446: begin cos_tmp = 24'b001010010001101010101011 ; sin_tmp = 24'b001100010000111000111001 ; end 
      12'd447: begin cos_tmp = 24'b001010001111001100101010 ; sin_tmp = 24'b001100010010111100111000 ; end 
      12'd448: begin cos_tmp = 24'b001010001111001100101010 ; sin_tmp = 24'b001100010010111100111000 ; end 
      12'd449: begin cos_tmp = 24'b001010001100101110001110 ; sin_tmp = 24'b001100010101000000010111 ; end 
      12'd450: begin cos_tmp = 24'b001010001010001111011000 ; sin_tmp = 24'b001100010111000011010110 ; end 
      12'd451: begin cos_tmp = 24'b001010001010001111011000 ; sin_tmp = 24'b001100010111000011010110 ; end 
      12'd452: begin cos_tmp = 24'b001010000111110000001000 ; sin_tmp = 24'b001100011001000101110101 ; end 
      12'd453: begin cos_tmp = 24'b001010000111110000001000 ; sin_tmp = 24'b001100011001000101110101 ; end 
      12'd454: begin cos_tmp = 24'b001010000101010000011101 ; sin_tmp = 24'b001100011011000111110100 ; end 
      12'd455: begin cos_tmp = 24'b001010000010110000011000 ; sin_tmp = 24'b001100011101001001010100 ; end 
      12'd456: begin cos_tmp = 24'b001010000010110000011000 ; sin_tmp = 24'b001100011101001001010100 ; end 
      12'd457: begin cos_tmp = 24'b001010000000001111111010 ; sin_tmp = 24'b001100011111001010010010 ; end 
      12'd458: begin cos_tmp = 24'b001001111101101111000001 ; sin_tmp = 24'b001100100001001010110001 ; end 
      12'd459: begin cos_tmp = 24'b001001111101101111000001 ; sin_tmp = 24'b001100100001001010110001 ; end 
      12'd460: begin cos_tmp = 24'b001001111011001101101111 ; sin_tmp = 24'b001100100011001010101111 ; end 
      12'd461: begin cos_tmp = 24'b001001111011001101101111 ; sin_tmp = 24'b001100100011001010101111 ; end 
      12'd462: begin cos_tmp = 24'b001001111000101100000011 ; sin_tmp = 24'b001100100101001010001101 ; end 
      12'd463: begin cos_tmp = 24'b001001110110001001111110 ; sin_tmp = 24'b001100100111001001001010 ; end 
      12'd464: begin cos_tmp = 24'b001001110110001001111110 ; sin_tmp = 24'b001100100111001001001010 ; end 
      12'd465: begin cos_tmp = 24'b001001110011100111011111 ; sin_tmp = 24'b001100101001000111100110 ; end 
      12'd466: begin cos_tmp = 24'b001001110001000100100110 ; sin_tmp = 24'b001100101011000101100010 ; end 
      12'd467: begin cos_tmp = 24'b001001110001000100100110 ; sin_tmp = 24'b001100101011000101100010 ; end 
      12'd468: begin cos_tmp = 24'b001001101110100001010100 ; sin_tmp = 24'b001100101101000010111101 ; end 
      12'd469: begin cos_tmp = 24'b001001101110100001010100 ; sin_tmp = 24'b001100101101000010111101 ; end 
      12'd470: begin cos_tmp = 24'b001001101011111101101010 ; sin_tmp = 24'b001100101110111111110111 ; end 
      12'd471: begin cos_tmp = 24'b001001101001011001100110 ; sin_tmp = 24'b001100110000111100010000 ; end 
      12'd472: begin cos_tmp = 24'b001001101001011001100110 ; sin_tmp = 24'b001100110000111100010000 ; end 
      12'd473: begin cos_tmp = 24'b001001100110110101001001 ; sin_tmp = 24'b001100110010111000001001 ; end 
      12'd474: begin cos_tmp = 24'b001001100110110101001001 ; sin_tmp = 24'b001100110010111000001001 ; end 
      12'd475: begin cos_tmp = 24'b001001100100010000010011 ; sin_tmp = 24'b001100110100110011100000 ; end 
      12'd476: begin cos_tmp = 24'b001001100001101011000101 ; sin_tmp = 24'b001100110110101110010101 ; end 
      12'd477: begin cos_tmp = 24'b001001100001101011000101 ; sin_tmp = 24'b001100110110101110010101 ; end 
      12'd478: begin cos_tmp = 24'b001001011111000101011110 ; sin_tmp = 24'b001100111000101000101010 ; end 
      12'd479: begin cos_tmp = 24'b001001011100011111011110 ; sin_tmp = 24'b001100111010100010011101 ; end 
      12'd480: begin cos_tmp = 24'b001001011100011111011110 ; sin_tmp = 24'b001100111010100010011101 ; end 
      12'd481: begin cos_tmp = 24'b001001011001111001000110 ; sin_tmp = 24'b001100111100011011101111 ; end 
      12'd482: begin cos_tmp = 24'b001001011001111001000110 ; sin_tmp = 24'b001100111100011011101111 ; end 
      12'd483: begin cos_tmp = 24'b001001010111010010010110 ; sin_tmp = 24'b001100111110010100100000 ; end 
      12'd484: begin cos_tmp = 24'b001001010100101011001101 ; sin_tmp = 24'b001101000000001100101110 ; end 
      12'd485: begin cos_tmp = 24'b001001010100101011001101 ; sin_tmp = 24'b001101000000001100101110 ; end 
      12'd486: begin cos_tmp = 24'b001001010010000011101100 ; sin_tmp = 24'b001101000010000100011100 ; end 
      12'd487: begin cos_tmp = 24'b001001001111011011110100 ; sin_tmp = 24'b001101000011111011100111 ; end 
      12'd488: begin cos_tmp = 24'b001001001111011011110100 ; sin_tmp = 24'b001101000011111011100111 ; end 
      12'd489: begin cos_tmp = 24'b001001001100110011100011 ; sin_tmp = 24'b001101000101110010010001 ; end 
      12'd490: begin cos_tmp = 24'b001001001100110011100011 ; sin_tmp = 24'b001101000101110010010001 ; end 
      12'd491: begin cos_tmp = 24'b001001001010001010111010 ; sin_tmp = 24'b001101000111101000011000 ; end 
      12'd492: begin cos_tmp = 24'b001001000111100001111010 ; sin_tmp = 24'b001101001001011101111110 ; end 
      12'd493: begin cos_tmp = 24'b001001000111100001111010 ; sin_tmp = 24'b001101001001011101111110 ; end 
      12'd494: begin cos_tmp = 24'b001001000100111000100010 ; sin_tmp = 24'b001101001011010011000010 ; end 
      12'd495: begin cos_tmp = 24'b001001000010001110110011 ; sin_tmp = 24'b001101001101000111100100 ; end 
      12'd496: begin cos_tmp = 24'b001001000010001110110011 ; sin_tmp = 24'b001101001101000111100100 ; end 
      12'd497: begin cos_tmp = 24'b001000111111100100101101 ; sin_tmp = 24'b001101001110111011100011 ; end 
      12'd498: begin cos_tmp = 24'b001000111111100100101101 ; sin_tmp = 24'b001101001110111011100011 ; end 
      12'd499: begin cos_tmp = 24'b001000111100111010001111 ; sin_tmp = 24'b001101010000101111000001 ; end 
      12'd500: begin cos_tmp = 24'b001000111010001111011010 ; sin_tmp = 24'b001101010010100001111100 ; end 
      12'd501: begin cos_tmp = 24'b001000111010001111011010 ; sin_tmp = 24'b001101010010100001111100 ; end 
      12'd502: begin cos_tmp = 24'b001000110111100100001110 ; sin_tmp = 24'b001101010100010100010100 ; end 
      12'd503: begin cos_tmp = 24'b001000110100111000101010 ; sin_tmp = 24'b001101010110000110001011 ; end 
      12'd504: begin cos_tmp = 24'b001000110100111000101010 ; sin_tmp = 24'b001101010110000110001011 ; end 
      12'd505: begin cos_tmp = 24'b001000110010001100110001 ; sin_tmp = 24'b001101010111110111011110 ; end 
      12'd506: begin cos_tmp = 24'b001000110010001100110001 ; sin_tmp = 24'b001101010111110111011110 ; end 
      12'd507: begin cos_tmp = 24'b001000101111100000100000 ; sin_tmp = 24'b001101011001101000001111 ; end 
      12'd508: begin cos_tmp = 24'b001000101100110011111001 ; sin_tmp = 24'b001101011011011000011110 ; end 
      12'd509: begin cos_tmp = 24'b001000101100110011111001 ; sin_tmp = 24'b001101011011011000011110 ; end 
      12'd510: begin cos_tmp = 24'b001000101010000110111011 ; sin_tmp = 24'b001101011101001000001001 ; end 
      12'd511: begin cos_tmp = 24'b001000101010000110111011 ; sin_tmp = 24'b001101011101001000001001 ; end 
      12'd512: begin cos_tmp = 24'b001000100111011001100111 ; sin_tmp = 24'b001101011110110111010010 ; end 
      12'd513: begin cos_tmp = 24'b001000100100101011111100 ; sin_tmp = 24'b001101100000100101111000 ; end 
      12'd514: begin cos_tmp = 24'b001000100100101011111100 ; sin_tmp = 24'b001101100000100101111000 ; end 
      12'd515: begin cos_tmp = 24'b001000100001111101111100 ; sin_tmp = 24'b001101100010010011111011 ; end 
      12'd516: begin cos_tmp = 24'b001000011111001111100101 ; sin_tmp = 24'b001101100100000001011011 ; end 
      12'd517: begin cos_tmp = 24'b001000011111001111100101 ; sin_tmp = 24'b001101100100000001011011 ; end 
      12'd518: begin cos_tmp = 24'b001000011100100000111001 ; sin_tmp = 24'b001101100101101110011000 ; end 
      12'd519: begin cos_tmp = 24'b001000011100100000111001 ; sin_tmp = 24'b001101100101101110011000 ; end 
      12'd520: begin cos_tmp = 24'b001000011001110001110110 ; sin_tmp = 24'b001101100111011010110010 ; end 
      12'd521: begin cos_tmp = 24'b001000010111000010011110 ; sin_tmp = 24'b001101101001000110101000 ; end 
      12'd522: begin cos_tmp = 24'b001000010111000010011110 ; sin_tmp = 24'b001101101001000110101000 ; end 
      12'd523: begin cos_tmp = 24'b001000010100010010110000 ; sin_tmp = 24'b001101101010110001111011 ; end 
      12'd524: begin cos_tmp = 24'b001000010001100010101101 ; sin_tmp = 24'b001101101100011100101011 ; end 
      12'd525: begin cos_tmp = 24'b001000010001100010101101 ; sin_tmp = 24'b001101101100011100101011 ; end 
      12'd526: begin cos_tmp = 24'b001000001110110010010100 ; sin_tmp = 24'b001101101110000110110111 ; end 
      12'd527: begin cos_tmp = 24'b001000001110110010010100 ; sin_tmp = 24'b001101101110000110110111 ; end 
      12'd528: begin cos_tmp = 24'b001000001100000001100110 ; sin_tmp = 24'b001101101111110000100000 ; end 
      12'd529: begin cos_tmp = 24'b001000001001010000100010 ; sin_tmp = 24'b001101110001011001100110 ; end 
      12'd530: begin cos_tmp = 24'b001000001001010000100010 ; sin_tmp = 24'b001101110001011001100110 ; end 
      12'd531: begin cos_tmp = 24'b001000000110011111001010 ; sin_tmp = 24'b001101110011000010000111 ; end 
      12'd532: begin cos_tmp = 24'b001000000011101101011101 ; sin_tmp = 24'b001101110100101010000101 ; end 
      12'd533: begin cos_tmp = 24'b001000000011101101011101 ; sin_tmp = 24'b001101110100101010000101 ; end 
      12'd534: begin cos_tmp = 24'b001000000000111011011011 ; sin_tmp = 24'b001101110110010001100000 ; end 
      12'd535: begin cos_tmp = 24'b001000000000111011011011 ; sin_tmp = 24'b001101110110010001100000 ; end 
      12'd536: begin cos_tmp = 24'b000111111110001001000100 ; sin_tmp = 24'b001101110111111000010110 ; end 
      12'd537: begin cos_tmp = 24'b000111111011010110011000 ; sin_tmp = 24'b001101111001011110101001 ; end 
      12'd538: begin cos_tmp = 24'b000111111011010110011000 ; sin_tmp = 24'b001101111001011110101001 ; end 
      12'd539: begin cos_tmp = 24'b000111111000100011011000 ; sin_tmp = 24'b001101111011000100010111 ; end 
      12'd540: begin cos_tmp = 24'b000111110101110000000100 ; sin_tmp = 24'b001101111100101001100010 ; end 
      12'd541: begin cos_tmp = 24'b000111110101110000000100 ; sin_tmp = 24'b001101111100101001100010 ; end 
      12'd542: begin cos_tmp = 24'b000111110010111100011011 ; sin_tmp = 24'b001101111110001110001000 ; end 
      12'd543: begin cos_tmp = 24'b000111110010111100011011 ; sin_tmp = 24'b001101111110001110001000 ; end 
      12'd544: begin cos_tmp = 24'b000111110000001000011110 ; sin_tmp = 24'b001101111111110010001011 ; end 
      12'd545: begin cos_tmp = 24'b000111101101010100001101 ; sin_tmp = 24'b001110000001010101101001 ; end 
      12'd546: begin cos_tmp = 24'b000111101101010100001101 ; sin_tmp = 24'b001110000001010101101001 ; end 
      12'd547: begin cos_tmp = 24'b000111101010011111101000 ; sin_tmp = 24'b001110000010111000100010 ; end 
      12'd548: begin cos_tmp = 24'b000111100111101010110000 ; sin_tmp = 24'b001110000100011010111000 ; end 
      12'd549: begin cos_tmp = 24'b000111100111101010110000 ; sin_tmp = 24'b001110000100011010111000 ; end 
      12'd550: begin cos_tmp = 24'b000111100100110101100011 ; sin_tmp = 24'b001110000101111100101001 ; end 
      12'd551: begin cos_tmp = 24'b000111100100110101100011 ; sin_tmp = 24'b001110000101111100101001 ; end 
      12'd552: begin cos_tmp = 24'b000111100010000000000011 ; sin_tmp = 24'b001110000111011101110110 ; end 
      12'd553: begin cos_tmp = 24'b000111011111001010010000 ; sin_tmp = 24'b001110001000111110011110 ; end 
      12'd554: begin cos_tmp = 24'b000111011111001010010000 ; sin_tmp = 24'b001110001000111110011110 ; end 
      12'd555: begin cos_tmp = 24'b000111011100010100001001 ; sin_tmp = 24'b001110001010011110100001 ; end 
      12'd556: begin cos_tmp = 24'b000111011100010100001001 ; sin_tmp = 24'b001110001010011110100001 ; end 
      12'd557: begin cos_tmp = 24'b000111011001011101101111 ; sin_tmp = 24'b001110001011111110000000 ; end 
      12'd558: begin cos_tmp = 24'b000111010110100111000010 ; sin_tmp = 24'b001110001101011100111010 ; end 
      12'd559: begin cos_tmp = 24'b000111010110100111000010 ; sin_tmp = 24'b001110001101011100111010 ; end 
      12'd560: begin cos_tmp = 24'b000111010011110000000001 ; sin_tmp = 24'b001110001110111011010000 ; end 
      12'd561: begin cos_tmp = 24'b000111010000111000101110 ; sin_tmp = 24'b001110010000011001000000 ; end 
      12'd562: begin cos_tmp = 24'b000111010000111000101110 ; sin_tmp = 24'b001110010000011001000000 ; end 
      12'd563: begin cos_tmp = 24'b000111001110000001001000 ; sin_tmp = 24'b001110010001110110001100 ; end 
      12'd564: begin cos_tmp = 24'b000111001110000001001000 ; sin_tmp = 24'b001110010001110110001100 ; end 
      12'd565: begin cos_tmp = 24'b000111001011001001010000 ; sin_tmp = 24'b001110010011010010110011 ; end 
      12'd566: begin cos_tmp = 24'b000111001000010001000100 ; sin_tmp = 24'b001110010100101110110100 ; end 
      12'd567: begin cos_tmp = 24'b000111001000010001000100 ; sin_tmp = 24'b001110010100101110110100 ; end 
      12'd568: begin cos_tmp = 24'b000111000101011000100111 ; sin_tmp = 24'b001110010110001010010001 ; end 
      12'd569: begin cos_tmp = 24'b000111000010011111110111 ; sin_tmp = 24'b001110010111100101001001 ; end 
      12'd570: begin cos_tmp = 24'b000111000010011111110111 ; sin_tmp = 24'b001110010111100101001001 ; end 
      12'd571: begin cos_tmp = 24'b000110111111100110110100 ; sin_tmp = 24'b001110011000111111011011 ; end 
      12'd572: begin cos_tmp = 24'b000110111111100110110100 ; sin_tmp = 24'b001110011000111111011011 ; end 
      12'd573: begin cos_tmp = 24'b000110111100101101100000 ; sin_tmp = 24'b001110011010011001001000 ; end 
      12'd574: begin cos_tmp = 24'b000110111001110011111010 ; sin_tmp = 24'b001110011011110010010000 ; end 
      12'd575: begin cos_tmp = 24'b000110111001110011111010 ; sin_tmp = 24'b001110011011110010010000 ; end 
      12'd576: begin cos_tmp = 24'b000110110110111010000010 ; sin_tmp = 24'b001110011101001010110011 ; end 
      12'd577: begin cos_tmp = 24'b000110110011111111111000 ; sin_tmp = 24'b001110011110100010110000 ; end 
      12'd578: begin cos_tmp = 24'b000110110011111111111000 ; sin_tmp = 24'b001110011110100010110000 ; end 
      12'd579: begin cos_tmp = 24'b000110110001000101011100 ; sin_tmp = 24'b001110011111111010000111 ; end 
      12'd580: begin cos_tmp = 24'b000110110001000101011100 ; sin_tmp = 24'b001110011111111010000111 ; end 
      12'd581: begin cos_tmp = 24'b000110101110001010101111 ; sin_tmp = 24'b001110100001010000111010 ; end 
      12'd582: begin cos_tmp = 24'b000110101011001111110001 ; sin_tmp = 24'b001110100010100111000110 ; end 
      12'd583: begin cos_tmp = 24'b000110101011001111110001 ; sin_tmp = 24'b001110100010100111000110 ; end 
      12'd584: begin cos_tmp = 24'b000110101000010100100001 ; sin_tmp = 24'b001110100011111100101101 ; end 
      12'd585: begin cos_tmp = 24'b000110100101011001000000 ; sin_tmp = 24'b001110100101010001101110 ; end 
      12'd586: begin cos_tmp = 24'b000110100101011001000000 ; sin_tmp = 24'b001110100101010001101110 ; end 
      12'd587: begin cos_tmp = 24'b000110100010011101001110 ; sin_tmp = 24'b001110100110100110001010 ; end 
      12'd588: begin cos_tmp = 24'b000110100010011101001110 ; sin_tmp = 24'b001110100110100110001010 ; end 
      12'd589: begin cos_tmp = 24'b000110011111100001001100 ; sin_tmp = 24'b001110100111111010000000 ; end 
      12'd590: begin cos_tmp = 24'b000110011100100100111000 ; sin_tmp = 24'b001110101001001101010000 ; end 
      12'd591: begin cos_tmp = 24'b000110011100100100111000 ; sin_tmp = 24'b001110101001001101010000 ; end 
      12'd592: begin cos_tmp = 24'b000110011001101000010100 ; sin_tmp = 24'b001110101010011111111010 ; end 
      12'd593: begin cos_tmp = 24'b000110011001101000010100 ; sin_tmp = 24'b001110101010011111111010 ; end 
      12'd594: begin cos_tmp = 24'b000110010110101011011111 ; sin_tmp = 24'b001110101011110001111110 ; end 
      12'd595: begin cos_tmp = 24'b000110010011101110011010 ; sin_tmp = 24'b001110101101000011011100 ; end 
      12'd596: begin cos_tmp = 24'b000110010011101110011010 ; sin_tmp = 24'b001110101101000011011100 ; end 
      12'd597: begin cos_tmp = 24'b000110010000110001000100 ; sin_tmp = 24'b001110101110010100010100 ; end 
      12'd598: begin cos_tmp = 24'b000110001101110011011110 ; sin_tmp = 24'b001110101111100100100110 ; end 
      12'd599: begin cos_tmp = 24'b000110001101110011011110 ; sin_tmp = 24'b001110101111100100100110 ; end 
      12'd600: begin cos_tmp = 24'b000110001010110101101000 ; sin_tmp = 24'b001110110000110100010010 ; end 
      12'd601: begin cos_tmp = 24'b000110001010110101101000 ; sin_tmp = 24'b001110110000110100010010 ; end 
      12'd602: begin cos_tmp = 24'b000110000111110111100011 ; sin_tmp = 24'b001110110010000011011000 ; end 
      12'd603: begin cos_tmp = 24'b000110000100111001001101 ; sin_tmp = 24'b001110110011010001110111 ; end 
      12'd604: begin cos_tmp = 24'b000110000100111001001101 ; sin_tmp = 24'b001110110011010001110111 ; end 
      12'd605: begin cos_tmp = 24'b000110000001111010101000 ; sin_tmp = 24'b001110110100011111110000 ; end 
      12'd606: begin cos_tmp = 24'b000101111110111011110011 ; sin_tmp = 24'b001110110101101101000011 ; end 
      12'd607: begin cos_tmp = 24'b000101111110111011110011 ; sin_tmp = 24'b001110110101101101000011 ; end 
      12'd608: begin cos_tmp = 24'b000101111011111100101110 ; sin_tmp = 24'b001110110110111001101111 ; end 
      12'd609: begin cos_tmp = 24'b000101111011111100101110 ; sin_tmp = 24'b001110110110111001101111 ; end 
      12'd610: begin cos_tmp = 24'b000101111000111101011010 ; sin_tmp = 24'b001110111000000101110101 ; end 
      12'd611: begin cos_tmp = 24'b000101110101111101110111 ; sin_tmp = 24'b001110111001010001010101 ; end 
      12'd612: begin cos_tmp = 24'b000101110101111101110111 ; sin_tmp = 24'b001110111001010001010101 ; end 
      12'd613: begin cos_tmp = 24'b000101110010111110000101 ; sin_tmp = 24'b001110111010011100001110 ; end 
      12'd614: begin cos_tmp = 24'b000101101111111110000100 ; sin_tmp = 24'b001110111011100110100000 ; end 
      12'd615: begin cos_tmp = 24'b000101101111111110000100 ; sin_tmp = 24'b001110111011100110100000 ; end 
      12'd616: begin cos_tmp = 24'b000101101100111101110100 ; sin_tmp = 24'b001110111100110000001100 ; end 
      12'd617: begin cos_tmp = 24'b000101101100111101110100 ; sin_tmp = 24'b001110111100110000001100 ; end 
      12'd618: begin cos_tmp = 24'b000101101001111101010101 ; sin_tmp = 24'b001110111101111001010001 ; end 
      12'd619: begin cos_tmp = 24'b000101100110111100101000 ; sin_tmp = 24'b001110111111000001101111 ; end 
      12'd620: begin cos_tmp = 24'b000101100110111100101000 ; sin_tmp = 24'b001110111111000001101111 ; end 
      12'd621: begin cos_tmp = 24'b000101100011111011101100 ; sin_tmp = 24'b001111000000001001100110 ; end 
      12'd622: begin cos_tmp = 24'b000101100000111010100001 ; sin_tmp = 24'b001111000001010000110111 ; end 
      12'd623: begin cos_tmp = 24'b000101100000111010100001 ; sin_tmp = 24'b001111000001010000110111 ; end 
      12'd624: begin cos_tmp = 24'b000101011101111001001001 ; sin_tmp = 24'b001111000010010111100001 ; end 
      12'd625: begin cos_tmp = 24'b000101011101111001001001 ; sin_tmp = 24'b001111000010010111100001 ; end 
      12'd626: begin cos_tmp = 24'b000101011010110111100010 ; sin_tmp = 24'b001111000011011101100100 ; end 
      12'd627: begin cos_tmp = 24'b000101010111110101101101 ; sin_tmp = 24'b001111000100100011000000 ; end 
      12'd628: begin cos_tmp = 24'b000101010111110101101101 ; sin_tmp = 24'b001111000100100011000000 ; end 
      12'd629: begin cos_tmp = 24'b000101010100110011101010 ; sin_tmp = 24'b001111000101100111110101 ; end 
      12'd630: begin cos_tmp = 24'b000101010100110011101010 ; sin_tmp = 24'b001111000101100111110101 ; end 
      12'd631: begin cos_tmp = 24'b000101010001110001011010 ; sin_tmp = 24'b001111000110101100000011 ; end 
      12'd632: begin cos_tmp = 24'b000101001110101110111100 ; sin_tmp = 24'b001111000111101111101010 ; end 
      12'd633: begin cos_tmp = 24'b000101001110101110111100 ; sin_tmp = 24'b001111000111101111101010 ; end 
      12'd634: begin cos_tmp = 24'b000101001011101100010000 ; sin_tmp = 24'b001111001000110010101010 ; end 
      12'd635: begin cos_tmp = 24'b000101001000101001010111 ; sin_tmp = 24'b001111001001110101000010 ; end 
      12'd636: begin cos_tmp = 24'b000101001000101001010111 ; sin_tmp = 24'b001111001001110101000010 ; end 
      12'd637: begin cos_tmp = 24'b000101000101100110010001 ; sin_tmp = 24'b001111001010110110110100 ; end 
      12'd638: begin cos_tmp = 24'b000101000101100110010001 ; sin_tmp = 24'b001111001010110110110100 ; end 
      12'd639: begin cos_tmp = 24'b000101000010100010111101 ; sin_tmp = 24'b001111001011110111111110 ; end 
      12'd640: begin cos_tmp = 24'b000100111111011111011101 ; sin_tmp = 24'b001111001100111000100001 ; end 
      12'd641: begin cos_tmp = 24'b000100111111011111011101 ; sin_tmp = 24'b001111001100111000100001 ; end 
      12'd642: begin cos_tmp = 24'b000100111100011011101111 ; sin_tmp = 24'b001111001101111000011100 ; end 
      12'd643: begin cos_tmp = 24'b000100111001010111110101 ; sin_tmp = 24'b001111001110110111110000 ; end 
      12'd644: begin cos_tmp = 24'b000100111001010111110101 ; sin_tmp = 24'b001111001110110111110000 ; end 
      12'd645: begin cos_tmp = 24'b000100110110010011101110 ; sin_tmp = 24'b001111001111110110011101 ; end 
      12'd646: begin cos_tmp = 24'b000100110110010011101110 ; sin_tmp = 24'b001111001111110110011101 ; end 
      12'd647: begin cos_tmp = 24'b000100110011001111011011 ; sin_tmp = 24'b001111010000110100100010 ; end 
      12'd648: begin cos_tmp = 24'b000100110000001010111011 ; sin_tmp = 24'b001111010001110010000000 ; end 
      12'd649: begin cos_tmp = 24'b000100110000001010111011 ; sin_tmp = 24'b001111010001110010000000 ; end 
      12'd650: begin cos_tmp = 24'b000100101101000110001111 ; sin_tmp = 24'b001111010010101110110110 ; end 
      12'd651: begin cos_tmp = 24'b000100101010000001010110 ; sin_tmp = 24'b001111010011101011000101 ; end 
      12'd652: begin cos_tmp = 24'b000100101010000001010110 ; sin_tmp = 24'b001111010011101011000101 ; end 
      12'd653: begin cos_tmp = 24'b000100100110111100010010 ; sin_tmp = 24'b001111010100100110101100 ; end 
      12'd654: begin cos_tmp = 24'b000100100110111100010010 ; sin_tmp = 24'b001111010100100110101100 ; end 
      12'd655: begin cos_tmp = 24'b000100100011110111000001 ; sin_tmp = 24'b001111010101100001101100 ; end 
      12'd656: begin cos_tmp = 24'b000100100000110001100101 ; sin_tmp = 24'b001111010110011100000100 ; end 
      12'd657: begin cos_tmp = 24'b000100100000110001100101 ; sin_tmp = 24'b001111010110011100000100 ; end 
      12'd658: begin cos_tmp = 24'b000100011101101011111110 ; sin_tmp = 24'b001111010111010101110100 ; end 
      12'd659: begin cos_tmp = 24'b000100011010100110001010 ; sin_tmp = 24'b001111011000001110111100 ; end 
      12'd660: begin cos_tmp = 24'b000100011010100110001010 ; sin_tmp = 24'b001111011000001110111100 ; end 
      12'd661: begin cos_tmp = 24'b000100010111100000001011 ; sin_tmp = 24'b001111011001000111011101 ; end 
      12'd662: begin cos_tmp = 24'b000100010111100000001011 ; sin_tmp = 24'b001111011001000111011101 ; end 
      12'd663: begin cos_tmp = 24'b000100010100011010000001 ; sin_tmp = 24'b001111011001111111010101 ; end 
      12'd664: begin cos_tmp = 24'b000100010001010011101100 ; sin_tmp = 24'b001111011010110110100110 ; end 
      12'd665: begin cos_tmp = 24'b000100010001010011101100 ; sin_tmp = 24'b001111011010110110100110 ; end 
      12'd666: begin cos_tmp = 24'b000100001110001101001100 ; sin_tmp = 24'b001111011011101101001111 ; end 
      12'd667: begin cos_tmp = 24'b000100001110001101001100 ; sin_tmp = 24'b001111011011101101001111 ; end 
      12'd668: begin cos_tmp = 24'b000100001011000110100001 ; sin_tmp = 24'b001111011100100011010000 ; end 
      12'd669: begin cos_tmp = 24'b000100000111111111101011 ; sin_tmp = 24'b001111011101011000101001 ; end 
      12'd670: begin cos_tmp = 24'b000100000111111111101011 ; sin_tmp = 24'b001111011101011000101001 ; end 
      12'd671: begin cos_tmp = 24'b000100000100111000101010 ; sin_tmp = 24'b001111011110001101011010 ; end 
      12'd672: begin cos_tmp = 24'b000100000001110001011111 ; sin_tmp = 24'b001111011111000001100011 ; end 
      12'd673: begin cos_tmp = 24'b000100000001110001011111 ; sin_tmp = 24'b001111011111000001100011 ; end 
      12'd674: begin cos_tmp = 24'b000011111110101010001001 ; sin_tmp = 24'b001111011111110101000100 ; end 
      12'd675: begin cos_tmp = 24'b000011111110101010001001 ; sin_tmp = 24'b001111011111110101000100 ; end 
      12'd676: begin cos_tmp = 24'b000011111011100010101001 ; sin_tmp = 24'b001111100000100111111101 ; end 
      12'd677: begin cos_tmp = 24'b000011111000011010111111 ; sin_tmp = 24'b001111100001011010001110 ; end 
      12'd678: begin cos_tmp = 24'b000011111000011010111111 ; sin_tmp = 24'b001111100001011010001110 ; end 
      12'd679: begin cos_tmp = 24'b000011110101010011001011 ; sin_tmp = 24'b001111100010001011110110 ; end 
      12'd680: begin cos_tmp = 24'b000011110010001011001101 ; sin_tmp = 24'b001111100010111100110111 ; end 
      12'd681: begin cos_tmp = 24'b000011110010001011001101 ; sin_tmp = 24'b001111100010111100110111 ; end 
      12'd682: begin cos_tmp = 24'b000011101111000011000101 ; sin_tmp = 24'b001111100011101101001111 ; end 
      12'd683: begin cos_tmp = 24'b000011101111000011000101 ; sin_tmp = 24'b001111100011101101001111 ; end 
      12'd684: begin cos_tmp = 24'b000011101011111010110011 ; sin_tmp = 24'b001111100100011100111111 ; end 
      12'd685: begin cos_tmp = 24'b000011101000110010011000 ; sin_tmp = 24'b001111100101001100000111 ; end 
      12'd686: begin cos_tmp = 24'b000011101000110010011000 ; sin_tmp = 24'b001111100101001100000111 ; end 
      12'd687: begin cos_tmp = 24'b000011100101101001110100 ; sin_tmp = 24'b001111100101111010100110 ; end 
      12'd688: begin cos_tmp = 24'b000011100010100001000110 ; sin_tmp = 24'b001111100110101000011101 ; end 
      12'd689: begin cos_tmp = 24'b000011100010100001000110 ; sin_tmp = 24'b001111100110101000011101 ; end 
      12'd690: begin cos_tmp = 24'b000011011111011000001111 ; sin_tmp = 24'b001111100111010101101100 ; end 
      12'd691: begin cos_tmp = 24'b000011011111011000001111 ; sin_tmp = 24'b001111100111010101101100 ; end 
      12'd692: begin cos_tmp = 24'b000011011100001111001111 ; sin_tmp = 24'b001111101000000010010010 ; end 
      12'd693: begin cos_tmp = 24'b000011011001000110000110 ; sin_tmp = 24'b001111101000101110010000 ; end 
      12'd694: begin cos_tmp = 24'b000011011001000110000110 ; sin_tmp = 24'b001111101000101110010000 ; end 
      12'd695: begin cos_tmp = 24'b000011010101111100110101 ; sin_tmp = 24'b001111101001011001100101 ; end 
      12'd696: begin cos_tmp = 24'b000011010010110011011010 ; sin_tmp = 24'b001111101010000100010010 ; end 
      12'd697: begin cos_tmp = 24'b000011010010110011011010 ; sin_tmp = 24'b001111101010000100010010 ; end 
      12'd698: begin cos_tmp = 24'b000011001111101001111000 ; sin_tmp = 24'b001111101010101110010110 ; end 
      12'd699: begin cos_tmp = 24'b000011001111101001111000 ; sin_tmp = 24'b001111101010101110010110 ; end 
      12'd700: begin cos_tmp = 24'b000011001100100000001100 ; sin_tmp = 24'b001111101011010111110010 ; end 
      12'd701: begin cos_tmp = 24'b000011001001010110011001 ; sin_tmp = 24'b001111101100000000100101 ; end 
      12'd702: begin cos_tmp = 24'b000011001001010110011001 ; sin_tmp = 24'b001111101100000000100101 ; end 
      12'd703: begin cos_tmp = 24'b000011000110001100011101 ; sin_tmp = 24'b001111101100101000110000 ; end 
      12'd704: begin cos_tmp = 24'b000011000110001100011101 ; sin_tmp = 24'b001111101100101000110000 ; end 
      12'd705: begin cos_tmp = 24'b000011000011000010011010 ; sin_tmp = 24'b001111101101010000010010 ; end 
      12'd706: begin cos_tmp = 24'b000010111111111000001110 ; sin_tmp = 24'b001111101101110111001011 ; end 
      12'd707: begin cos_tmp = 24'b000010111111111000001110 ; sin_tmp = 24'b001111101101110111001011 ; end 
      12'd708: begin cos_tmp = 24'b000010111100101101111011 ; sin_tmp = 24'b001111101110011101011100 ; end 
      12'd709: begin cos_tmp = 24'b000010111001100011100000 ; sin_tmp = 24'b001111101111000011000100 ; end 
      12'd710: begin cos_tmp = 24'b000010111001100011100000 ; sin_tmp = 24'b001111101111000011000100 ; end 
      12'd711: begin cos_tmp = 24'b000010110110011000111110 ; sin_tmp = 24'b001111101111101000000100 ; end 
      12'd712: begin cos_tmp = 24'b000010110110011000111110 ; sin_tmp = 24'b001111101111101000000100 ; end 
      12'd713: begin cos_tmp = 24'b000010110011001110010100 ; sin_tmp = 24'b001111110000001100011010 ; end 
      12'd714: begin cos_tmp = 24'b000010110000000011100011 ; sin_tmp = 24'b001111110000110000001000 ; end 
      12'd715: begin cos_tmp = 24'b000010110000000011100011 ; sin_tmp = 24'b001111110000110000001000 ; end 
      12'd716: begin cos_tmp = 24'b000010101100111000101011 ; sin_tmp = 24'b001111110001010011001101 ; end 
      12'd717: begin cos_tmp = 24'b000010101001101101101100 ; sin_tmp = 24'b001111110001110101101001 ; end 
      12'd718: begin cos_tmp = 24'b000010101001101101101100 ; sin_tmp = 24'b001111110001110101101001 ; end 
      12'd719: begin cos_tmp = 24'b000010100110100010100110 ; sin_tmp = 24'b001111110010010111011101 ; end 
      12'd720: begin cos_tmp = 24'b000010100110100010100110 ; sin_tmp = 24'b001111110010010111011101 ; end 
      12'd721: begin cos_tmp = 24'b000010100011010111011001 ; sin_tmp = 24'b001111110010111000100111 ; end 
      12'd722: begin cos_tmp = 24'b000010100000001100000110 ; sin_tmp = 24'b001111110011011001001001 ; end 
      12'd723: begin cos_tmp = 24'b000010100000001100000110 ; sin_tmp = 24'b001111110011011001001001 ; end 
      12'd724: begin cos_tmp = 24'b000010011101000000101100 ; sin_tmp = 24'b001111110011111001000010 ; end 
      12'd725: begin cos_tmp = 24'b000010011001110101001100 ; sin_tmp = 24'b001111110100011000010010 ; end 
      12'd726: begin cos_tmp = 24'b000010011001110101001100 ; sin_tmp = 24'b001111110100011000010010 ; end 
      12'd727: begin cos_tmp = 24'b000010010110101001100101 ; sin_tmp = 24'b001111110100110110111001 ; end 
      12'd728: begin cos_tmp = 24'b000010010110101001100101 ; sin_tmp = 24'b001111110100110110111001 ; end 
      12'd729: begin cos_tmp = 24'b000010010011011101111001 ; sin_tmp = 24'b001111110101010100110111 ; end 
      12'd730: begin cos_tmp = 24'b000010010000010010000111 ; sin_tmp = 24'b001111110101110010001100 ; end 
      12'd731: begin cos_tmp = 24'b000010010000010010000111 ; sin_tmp = 24'b001111110101110010001100 ; end 
      12'd732: begin cos_tmp = 24'b000010001101000110001110 ; sin_tmp = 24'b001111110110001110111000 ; end 
      12'd733: begin cos_tmp = 24'b000010001001111010010000 ; sin_tmp = 24'b001111110110101010111011 ; end 
      12'd734: begin cos_tmp = 24'b000010001001111010010000 ; sin_tmp = 24'b001111110110101010111011 ; end 
      12'd735: begin cos_tmp = 24'b000010000110101110001101 ; sin_tmp = 24'b001111110111000110010110 ; end 
      12'd736: begin cos_tmp = 24'b000010000110101110001101 ; sin_tmp = 24'b001111110111000110010110 ; end 
      12'd737: begin cos_tmp = 24'b000010000011100010000100 ; sin_tmp = 24'b001111110111100001000111 ; end 
      12'd738: begin cos_tmp = 24'b000010000000010101110110 ; sin_tmp = 24'b001111110111111011001111 ; end 
      12'd739: begin cos_tmp = 24'b000010000000010101110110 ; sin_tmp = 24'b001111110111111011001111 ; end 
      12'd740: begin cos_tmp = 24'b000001111101001001100010 ; sin_tmp = 24'b001111111000010100101110 ; end 
      12'd741: begin cos_tmp = 24'b000001111101001001100010 ; sin_tmp = 24'b001111111000010100101110 ; end 
      12'd742: begin cos_tmp = 24'b000001111001111101001010 ; sin_tmp = 24'b001111111000101101100011 ; end 
      12'd743: begin cos_tmp = 24'b000001110110110000101100 ; sin_tmp = 24'b001111111001000101110000 ; end 
      12'd744: begin cos_tmp = 24'b000001110110110000101100 ; sin_tmp = 24'b001111111001000101110000 ; end 
      12'd745: begin cos_tmp = 24'b000001110011100100001010 ; sin_tmp = 24'b001111111001011101010100 ; end 
      12'd746: begin cos_tmp = 24'b000001110000010111100011 ; sin_tmp = 24'b001111111001110100001110 ; end 
      12'd747: begin cos_tmp = 24'b000001110000010111100011 ; sin_tmp = 24'b001111111001110100001110 ; end 
      12'd748: begin cos_tmp = 24'b000001101101001010111000 ; sin_tmp = 24'b001111111010001010100000 ; end 
      12'd749: begin cos_tmp = 24'b000001101101001010111000 ; sin_tmp = 24'b001111111010001010100000 ; end 
      12'd750: begin cos_tmp = 24'b000001101001111110001000 ; sin_tmp = 24'b001111111010100000001000 ; end 
      12'd751: begin cos_tmp = 24'b000001100110110001010100 ; sin_tmp = 24'b001111111010110101000111 ; end 
      12'd752: begin cos_tmp = 24'b000001100110110001010100 ; sin_tmp = 24'b001111111010110101000111 ; end 
      12'd753: begin cos_tmp = 24'b000001100011100100011011 ; sin_tmp = 24'b001111111011001001011101 ; end 
      12'd754: begin cos_tmp = 24'b000001100000010111011111 ; sin_tmp = 24'b001111111011011101001010 ; end 
      12'd755: begin cos_tmp = 24'b000001100000010111011111 ; sin_tmp = 24'b001111111011011101001010 ; end 
      12'd756: begin cos_tmp = 24'b000001011101001010011111 ; sin_tmp = 24'b001111111011110000001101 ; end 
      12'd757: begin cos_tmp = 24'b000001011101001010011111 ; sin_tmp = 24'b001111111011110000001101 ; end 
      12'd758: begin cos_tmp = 24'b000001011001111101011011 ; sin_tmp = 24'b001111111100000010100111 ; end 
      12'd759: begin cos_tmp = 24'b000001010110110000010011 ; sin_tmp = 24'b001111111100010100011000 ; end 
      12'd760: begin cos_tmp = 24'b000001010110110000010011 ; sin_tmp = 24'b001111111100010100011000 ; end 
      12'd761: begin cos_tmp = 24'b000001010011100011001000 ; sin_tmp = 24'b001111111100100101100000 ; end 
      12'd762: begin cos_tmp = 24'b000001010000010101111001 ; sin_tmp = 24'b001111111100110101111110 ; end 
      12'd763: begin cos_tmp = 24'b000001010000010101111001 ; sin_tmp = 24'b001111111100110101111110 ; end 
      12'd764: begin cos_tmp = 24'b000001001101001000101000 ; sin_tmp = 24'b001111111101000101110100 ; end 
      12'd765: begin cos_tmp = 24'b000001001101001000101000 ; sin_tmp = 24'b001111111101000101110100 ; end 
      12'd766: begin cos_tmp = 24'b000001001001111011010011 ; sin_tmp = 24'b001111111101010100111111 ; end 
      12'd767: begin cos_tmp = 24'b000001000110101101111011 ; sin_tmp = 24'b001111111101100011100010 ; end 
      12'd768: begin cos_tmp = 24'b000001000110101101111011 ; sin_tmp = 24'b001111111101100011100010 ; end 
      12'd769: begin cos_tmp = 24'b000001000011100000100000 ; sin_tmp = 24'b001111111101110001011011 ; end 
      12'd770: begin cos_tmp = 24'b000001000000010011000011 ; sin_tmp = 24'b001111111101111110101011 ; end 
      12'd771: begin cos_tmp = 24'b000001000000010011000011 ; sin_tmp = 24'b001111111101111110101011 ; end 
      12'd772: begin cos_tmp = 24'b000000111101000101100010 ; sin_tmp = 24'b001111111110001011010010 ; end 
      12'd773: begin cos_tmp = 24'b000000111101000101100010 ; sin_tmp = 24'b001111111110001011010010 ; end 
      12'd774: begin cos_tmp = 24'b000000111001111000000000 ; sin_tmp = 24'b001111111110010111010000 ; end 
      12'd775: begin cos_tmp = 24'b000000110110101010011011 ; sin_tmp = 24'b001111111110100010100100 ; end 
      12'd776: begin cos_tmp = 24'b000000110110101010011011 ; sin_tmp = 24'b001111111110100010100100 ; end 
      12'd777: begin cos_tmp = 24'b000000110011011100110100 ; sin_tmp = 24'b001111111110101101001110 ; end 
      12'd778: begin cos_tmp = 24'b000000110011011100110100 ; sin_tmp = 24'b001111111110101101001110 ; end 
      12'd779: begin cos_tmp = 24'b000000110000001111001011 ; sin_tmp = 24'b001111111110110111010000 ; end 
      12'd780: begin cos_tmp = 24'b000000101101000001100000 ; sin_tmp = 24'b001111111111000000101000 ; end 
      12'd781: begin cos_tmp = 24'b000000101101000001100000 ; sin_tmp = 24'b001111111111000000101000 ; end 
      12'd782: begin cos_tmp = 24'b000000101001110011110011 ; sin_tmp = 24'b001111111111001001010111 ; end 
      12'd783: begin cos_tmp = 24'b000000100110100110000100 ; sin_tmp = 24'b001111111111010001011100 ; end 
      12'd784: begin cos_tmp = 24'b000000100110100110000100 ; sin_tmp = 24'b001111111111010001011100 ; end 
      12'd785: begin cos_tmp = 24'b000000100011011000010100 ; sin_tmp = 24'b001111111111011000111000 ; end 
      12'd786: begin cos_tmp = 24'b000000100011011000010100 ; sin_tmp = 24'b001111111111011000111000 ; end 
      12'd787: begin cos_tmp = 24'b000000100000001010100010 ; sin_tmp = 24'b001111111111011111101010 ; end 
      12'd788: begin cos_tmp = 24'b000000011100111100101111 ; sin_tmp = 24'b001111111111100101110100 ; end 
      12'd789: begin cos_tmp = 24'b000000011100111100101111 ; sin_tmp = 24'b001111111111100101110100 ; end 
      12'd790: begin cos_tmp = 24'b000000011001101110111011 ; sin_tmp = 24'b001111111111101011010011 ; end 
      12'd791: begin cos_tmp = 24'b000000010110100001000110 ; sin_tmp = 24'b001111111111110000001010 ; end 
      12'd792: begin cos_tmp = 24'b000000010110100001000110 ; sin_tmp = 24'b001111111111110000001010 ; end 
      12'd793: begin cos_tmp = 24'b000000010011010011010000 ; sin_tmp = 24'b001111111111110100010111 ; end 
      12'd794: begin cos_tmp = 24'b000000010011010011010000 ; sin_tmp = 24'b001111111111110100010111 ; end 
      12'd795: begin cos_tmp = 24'b000000010000000101011001 ; sin_tmp = 24'b001111111111110111111011 ; end 
      12'd796: begin cos_tmp = 24'b000000001100110111100010 ; sin_tmp = 24'b001111111111111010110101 ; end 
      12'd797: begin cos_tmp = 24'b000000001100110111100010 ; sin_tmp = 24'b001111111111111010110101 ; end 
      12'd798: begin cos_tmp = 24'b000000001001101001101010 ; sin_tmp = 24'b001111111111111101000110 ; end 
      12'd799: begin cos_tmp = 24'b000000000110011011110001 ; sin_tmp = 24'b001111111111111110101101 ; end 
      12'd800: begin cos_tmp = 24'b000000000110011011110001 ; sin_tmp = 24'b001111111111111110101101 ; end 
      12'd801: begin cos_tmp = 24'b000000000011001101111001 ; sin_tmp = 24'b001111111111111111101011 ; end 
      12'd802: begin cos_tmp = 24'b000000000011001101111001 ; sin_tmp = 24'b001111111111111111101011 ; end 
      12'd803: begin cos_tmp = 24'b000000000000000000000000 ; sin_tmp = 24'b010000000000000000000000 ; end 
      
      endcase
      end
endmodule
