`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/08/17 23:58:24
// Design Name: 
// Module Name: cossin_16
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module cossin_16(
input wire signed [24:1] rad,
output  wire signed [16:1] cos,
output  wire signed [16:1] sin
    );
wire [1:0] sig ;
wire signed [24:1] rad_abs;
wire signed [24:1] rad_abs_90;
reg signed [16:1] cos_tmp;
reg signed [16:1] sin_tmp;

assign sig = {rad[24],rad_abs[24:13] > 805};
assign rad_abs = sig[1] ? - rad : rad ;
assign rad_abs_90 = sig[0] ? 24'd6588397- rad_abs : rad_abs; 
assign cos = sig[0] ? - cos_tmp : cos_tmp  ;
assign sin = sig[1] ? - sin_tmp : sin_tmp  ;
always @(*) begin
  case(rad_abs[24:13])
  12'd0: begin cos_tmp = 16'b0100000000000000 ; sin_tmp = 16'b0000000000110011 ; end 
  12'd1: begin cos_tmp = 16'b0100000000000000 ; sin_tmp = 16'b0000000000110011 ; end 
  12'd2: begin cos_tmp = 16'b0100000000000000 ; sin_tmp = 16'b0000000001100111 ; end 
  12'd3: begin cos_tmp = 16'b0011111111111111 ; sin_tmp = 16'b0000000010011010 ; end 
  12'd4: begin cos_tmp = 16'b0011111111111111 ; sin_tmp = 16'b0000000010011010 ; end 
  12'd5: begin cos_tmp = 16'b0011111111111111 ; sin_tmp = 16'b0000000011001110 ; end 
  12'd6: begin cos_tmp = 16'b0011111111111110 ; sin_tmp = 16'b0000000100000001 ; end 
  12'd7: begin cos_tmp = 16'b0011111111111110 ; sin_tmp = 16'b0000000100000001 ; end 
  12'd8: begin cos_tmp = 16'b0011111111111101 ; sin_tmp = 16'b0000000100110101 ; end 
  12'd9: begin cos_tmp = 16'b0011111111111101 ; sin_tmp = 16'b0000000100110101 ; end 
  12'd10: begin cos_tmp = 16'b0011111111111100 ; sin_tmp = 16'b0000000101101000 ; end 
  12'd11: begin cos_tmp = 16'b0011111111111011 ; sin_tmp = 16'b0000000110011100 ; end 
  12'd12: begin cos_tmp = 16'b0011111111111011 ; sin_tmp = 16'b0000000110011100 ; end 
  12'd13: begin cos_tmp = 16'b0011111111111001 ; sin_tmp = 16'b0000000111001111 ; end 
  12'd14: begin cos_tmp = 16'b0011111111111000 ; sin_tmp = 16'b0000001000000011 ; end 
  12'd15: begin cos_tmp = 16'b0011111111111000 ; sin_tmp = 16'b0000001000000011 ; end 
  12'd16: begin cos_tmp = 16'b0011111111110110 ; sin_tmp = 16'b0000001000110110 ; end 
  12'd17: begin cos_tmp = 16'b0011111111110110 ; sin_tmp = 16'b0000001000110110 ; end 
  12'd18: begin cos_tmp = 16'b0011111111110100 ; sin_tmp = 16'b0000001001101010 ; end 
  12'd19: begin cos_tmp = 16'b0011111111110010 ; sin_tmp = 16'b0000001010011101 ; end 
  12'd20: begin cos_tmp = 16'b0011111111110010 ; sin_tmp = 16'b0000001010011101 ; end 
  12'd21: begin cos_tmp = 16'b0011111111110000 ; sin_tmp = 16'b0000001011010000 ; end 
  12'd22: begin cos_tmp = 16'b0011111111110000 ; sin_tmp = 16'b0000001011010000 ; end 
  12'd23: begin cos_tmp = 16'b0011111111101110 ; sin_tmp = 16'b0000001100000100 ; end 
  12'd24: begin cos_tmp = 16'b0011111111101011 ; sin_tmp = 16'b0000001100110111 ; end 
  12'd25: begin cos_tmp = 16'b0011111111101011 ; sin_tmp = 16'b0000001100110111 ; end 
  12'd26: begin cos_tmp = 16'b0011111111101001 ; sin_tmp = 16'b0000001101101011 ; end 
  12'd27: begin cos_tmp = 16'b0011111111100110 ; sin_tmp = 16'b0000001110011110 ; end 
  12'd28: begin cos_tmp = 16'b0011111111100110 ; sin_tmp = 16'b0000001110011110 ; end 
  12'd29: begin cos_tmp = 16'b0011111111100011 ; sin_tmp = 16'b0000001111010001 ; end 
  12'd30: begin cos_tmp = 16'b0011111111100011 ; sin_tmp = 16'b0000001111010001 ; end 
  12'd31: begin cos_tmp = 16'b0011111111100000 ; sin_tmp = 16'b0000010000000101 ; end 
  12'd32: begin cos_tmp = 16'b0011111111011100 ; sin_tmp = 16'b0000010000111000 ; end 
  12'd33: begin cos_tmp = 16'b0011111111011100 ; sin_tmp = 16'b0000010000111000 ; end 
  12'd34: begin cos_tmp = 16'b0011111111011001 ; sin_tmp = 16'b0000010001101011 ; end 
  12'd35: begin cos_tmp = 16'b0011111111010101 ; sin_tmp = 16'b0000010010011111 ; end 
  12'd36: begin cos_tmp = 16'b0011111111010101 ; sin_tmp = 16'b0000010010011111 ; end 
  12'd37: begin cos_tmp = 16'b0011111111010001 ; sin_tmp = 16'b0000010011010010 ; end 
  12'd38: begin cos_tmp = 16'b0011111111010001 ; sin_tmp = 16'b0000010011010010 ; end 
  12'd39: begin cos_tmp = 16'b0011111111001101 ; sin_tmp = 16'b0000010100000101 ; end 
  12'd40: begin cos_tmp = 16'b0011111111001001 ; sin_tmp = 16'b0000010100111001 ; end 
  12'd41: begin cos_tmp = 16'b0011111111001001 ; sin_tmp = 16'b0000010100111001 ; end 
  12'd42: begin cos_tmp = 16'b0011111111000101 ; sin_tmp = 16'b0000010101101100 ; end 
  12'd43: begin cos_tmp = 16'b0011111111000001 ; sin_tmp = 16'b0000010110011111 ; end 
  12'd44: begin cos_tmp = 16'b0011111111000001 ; sin_tmp = 16'b0000010110011111 ; end 
  12'd45: begin cos_tmp = 16'b0011111110111100 ; sin_tmp = 16'b0000010111010011 ; end 
  12'd46: begin cos_tmp = 16'b0011111110111100 ; sin_tmp = 16'b0000010111010011 ; end 
  12'd47: begin cos_tmp = 16'b0011111110110111 ; sin_tmp = 16'b0000011000000110 ; end 
  12'd48: begin cos_tmp = 16'b0011111110110010 ; sin_tmp = 16'b0000011000111001 ; end 
  12'd49: begin cos_tmp = 16'b0011111110110010 ; sin_tmp = 16'b0000011000111001 ; end 
  12'd50: begin cos_tmp = 16'b0011111110101101 ; sin_tmp = 16'b0000011001101100 ; end 
  12'd51: begin cos_tmp = 16'b0011111110101000 ; sin_tmp = 16'b0000011010100000 ; end 
  12'd52: begin cos_tmp = 16'b0011111110101000 ; sin_tmp = 16'b0000011010100000 ; end 
  12'd53: begin cos_tmp = 16'b0011111110100011 ; sin_tmp = 16'b0000011011010011 ; end 
  12'd54: begin cos_tmp = 16'b0011111110100011 ; sin_tmp = 16'b0000011011010011 ; end 
  12'd55: begin cos_tmp = 16'b0011111110011101 ; sin_tmp = 16'b0000011100000110 ; end 
  12'd56: begin cos_tmp = 16'b0011111110010111 ; sin_tmp = 16'b0000011100111001 ; end 
  12'd57: begin cos_tmp = 16'b0011111110010111 ; sin_tmp = 16'b0000011100111001 ; end 
  12'd58: begin cos_tmp = 16'b0011111110010001 ; sin_tmp = 16'b0000011101101100 ; end 
  12'd59: begin cos_tmp = 16'b0011111110010001 ; sin_tmp = 16'b0000011101101100 ; end 
  12'd60: begin cos_tmp = 16'b0011111110001011 ; sin_tmp = 16'b0000011110011111 ; end 
  12'd61: begin cos_tmp = 16'b0011111110000101 ; sin_tmp = 16'b0000011111010010 ; end 
  12'd62: begin cos_tmp = 16'b0011111110000101 ; sin_tmp = 16'b0000011111010010 ; end 
  12'd63: begin cos_tmp = 16'b0011111101111111 ; sin_tmp = 16'b0000100000000101 ; end 
  12'd64: begin cos_tmp = 16'b0011111101111000 ; sin_tmp = 16'b0000100000111001 ; end 
  12'd65: begin cos_tmp = 16'b0011111101111000 ; sin_tmp = 16'b0000100000111001 ; end 
  12'd66: begin cos_tmp = 16'b0011111101110010 ; sin_tmp = 16'b0000100001101100 ; end 
  12'd67: begin cos_tmp = 16'b0011111101110010 ; sin_tmp = 16'b0000100001101100 ; end 
  12'd68: begin cos_tmp = 16'b0011111101101011 ; sin_tmp = 16'b0000100010011111 ; end 
  12'd69: begin cos_tmp = 16'b0011111101100100 ; sin_tmp = 16'b0000100011010010 ; end 
  12'd70: begin cos_tmp = 16'b0011111101100100 ; sin_tmp = 16'b0000100011010010 ; end 
  12'd71: begin cos_tmp = 16'b0011111101011101 ; sin_tmp = 16'b0000100100000101 ; end 
  12'd72: begin cos_tmp = 16'b0011111101010101 ; sin_tmp = 16'b0000100100110111 ; end 
  12'd73: begin cos_tmp = 16'b0011111101010101 ; sin_tmp = 16'b0000100100110111 ; end 
  12'd74: begin cos_tmp = 16'b0011111101001110 ; sin_tmp = 16'b0000100101101010 ; end 
  12'd75: begin cos_tmp = 16'b0011111101001110 ; sin_tmp = 16'b0000100101101010 ; end 
  12'd76: begin cos_tmp = 16'b0011111101000110 ; sin_tmp = 16'b0000100110011101 ; end 
  12'd77: begin cos_tmp = 16'b0011111100111110 ; sin_tmp = 16'b0000100111010000 ; end 
  12'd78: begin cos_tmp = 16'b0011111100111110 ; sin_tmp = 16'b0000100111010000 ; end 
  12'd79: begin cos_tmp = 16'b0011111100110110 ; sin_tmp = 16'b0000101000000011 ; end 
  12'd80: begin cos_tmp = 16'b0011111100101110 ; sin_tmp = 16'b0000101000110110 ; end 
  12'd81: begin cos_tmp = 16'b0011111100101110 ; sin_tmp = 16'b0000101000110110 ; end 
  12'd82: begin cos_tmp = 16'b0011111100100110 ; sin_tmp = 16'b0000101001101001 ; end 
  12'd83: begin cos_tmp = 16'b0011111100100110 ; sin_tmp = 16'b0000101001101001 ; end 
  12'd84: begin cos_tmp = 16'b0011111100011101 ; sin_tmp = 16'b0000101010011011 ; end 
  12'd85: begin cos_tmp = 16'b0011111100010101 ; sin_tmp = 16'b0000101011001110 ; end 
  12'd86: begin cos_tmp = 16'b0011111100010101 ; sin_tmp = 16'b0000101011001110 ; end 
  12'd87: begin cos_tmp = 16'b0011111100001100 ; sin_tmp = 16'b0000101100000001 ; end 
  12'd88: begin cos_tmp = 16'b0011111100000011 ; sin_tmp = 16'b0000101100110100 ; end 
  12'd89: begin cos_tmp = 16'b0011111100000011 ; sin_tmp = 16'b0000101100110100 ; end 
  12'd90: begin cos_tmp = 16'b0011111011111010 ; sin_tmp = 16'b0000101101100110 ; end 
  12'd91: begin cos_tmp = 16'b0011111011111010 ; sin_tmp = 16'b0000101101100110 ; end 
  12'd92: begin cos_tmp = 16'b0011111011110001 ; sin_tmp = 16'b0000101110011001 ; end 
  12'd93: begin cos_tmp = 16'b0011111011100111 ; sin_tmp = 16'b0000101111001011 ; end 
  12'd94: begin cos_tmp = 16'b0011111011100111 ; sin_tmp = 16'b0000101111001011 ; end 
  12'd95: begin cos_tmp = 16'b0011111011011110 ; sin_tmp = 16'b0000101111111110 ; end 
  12'd96: begin cos_tmp = 16'b0011111011011110 ; sin_tmp = 16'b0000101111111110 ; end 
  12'd97: begin cos_tmp = 16'b0011111011010100 ; sin_tmp = 16'b0000110000110001 ; end 
  12'd98: begin cos_tmp = 16'b0011111011001010 ; sin_tmp = 16'b0000110001100011 ; end 
  12'd99: begin cos_tmp = 16'b0011111011001010 ; sin_tmp = 16'b0000110001100011 ; end 
  12'd100: begin cos_tmp = 16'b0011111011000000 ; sin_tmp = 16'b0000110010010110 ; end 
  12'd101: begin cos_tmp = 16'b0011111010110110 ; sin_tmp = 16'b0000110011001000 ; end 
  12'd102: begin cos_tmp = 16'b0011111010110110 ; sin_tmp = 16'b0000110011001000 ; end 
  12'd103: begin cos_tmp = 16'b0011111010101100 ; sin_tmp = 16'b0000110011111010 ; end 
  12'd104: begin cos_tmp = 16'b0011111010101100 ; sin_tmp = 16'b0000110011111010 ; end 
  12'd105: begin cos_tmp = 16'b0011111010100001 ; sin_tmp = 16'b0000110100101101 ; end 
  12'd106: begin cos_tmp = 16'b0011111010010110 ; sin_tmp = 16'b0000110101011111 ; end 
  12'd107: begin cos_tmp = 16'b0011111010010110 ; sin_tmp = 16'b0000110101011111 ; end 
  12'd108: begin cos_tmp = 16'b0011111010001100 ; sin_tmp = 16'b0000110110010010 ; end 
  12'd109: begin cos_tmp = 16'b0011111010000001 ; sin_tmp = 16'b0000110111000100 ; end 
  12'd110: begin cos_tmp = 16'b0011111010000001 ; sin_tmp = 16'b0000110111000100 ; end 
  12'd111: begin cos_tmp = 16'b0011111001110101 ; sin_tmp = 16'b0000110111110110 ; end 
  12'd112: begin cos_tmp = 16'b0011111001110101 ; sin_tmp = 16'b0000110111110110 ; end 
  12'd113: begin cos_tmp = 16'b0011111001101010 ; sin_tmp = 16'b0000111000101000 ; end 
  12'd114: begin cos_tmp = 16'b0011111001011111 ; sin_tmp = 16'b0000111001011010 ; end 
  12'd115: begin cos_tmp = 16'b0011111001011111 ; sin_tmp = 16'b0000111001011010 ; end 
  12'd116: begin cos_tmp = 16'b0011111001010011 ; sin_tmp = 16'b0000111010001101 ; end 
  12'd117: begin cos_tmp = 16'b0011111001000111 ; sin_tmp = 16'b0000111010111111 ; end 
  12'd118: begin cos_tmp = 16'b0011111001000111 ; sin_tmp = 16'b0000111010111111 ; end 
  12'd119: begin cos_tmp = 16'b0011111000111011 ; sin_tmp = 16'b0000111011110001 ; end 
  12'd120: begin cos_tmp = 16'b0011111000111011 ; sin_tmp = 16'b0000111011110001 ; end 
  12'd121: begin cos_tmp = 16'b0011111000101111 ; sin_tmp = 16'b0000111100100011 ; end 
  12'd122: begin cos_tmp = 16'b0011111000100011 ; sin_tmp = 16'b0000111101010101 ; end 
  12'd123: begin cos_tmp = 16'b0011111000100011 ; sin_tmp = 16'b0000111101010101 ; end 
  12'd124: begin cos_tmp = 16'b0011111000010111 ; sin_tmp = 16'b0000111110000111 ; end 
  12'd125: begin cos_tmp = 16'b0011111000001010 ; sin_tmp = 16'b0000111110111001 ; end 
  12'd126: begin cos_tmp = 16'b0011111000001010 ; sin_tmp = 16'b0000111110111001 ; end 
  12'd127: begin cos_tmp = 16'b0011110111111101 ; sin_tmp = 16'b0000111111101011 ; end 
  12'd128: begin cos_tmp = 16'b0011110111111101 ; sin_tmp = 16'b0000111111101011 ; end 
  12'd129: begin cos_tmp = 16'b0011110111110000 ; sin_tmp = 16'b0001000000011100 ; end 
  12'd130: begin cos_tmp = 16'b0011110111100011 ; sin_tmp = 16'b0001000001001110 ; end 
  12'd131: begin cos_tmp = 16'b0011110111100011 ; sin_tmp = 16'b0001000001001110 ; end 
  12'd132: begin cos_tmp = 16'b0011110111010110 ; sin_tmp = 16'b0001000010000000 ; end 
  12'd133: begin cos_tmp = 16'b0011110111010110 ; sin_tmp = 16'b0001000010000000 ; end 
  12'd134: begin cos_tmp = 16'b0011110111001001 ; sin_tmp = 16'b0001000010110010 ; end 
  12'd135: begin cos_tmp = 16'b0011110110111011 ; sin_tmp = 16'b0001000011100011 ; end 
  12'd136: begin cos_tmp = 16'b0011110110111011 ; sin_tmp = 16'b0001000011100011 ; end 
  12'd137: begin cos_tmp = 16'b0011110110101110 ; sin_tmp = 16'b0001000100010101 ; end 
  12'd138: begin cos_tmp = 16'b0011110110100000 ; sin_tmp = 16'b0001000101000111 ; end 
  12'd139: begin cos_tmp = 16'b0011110110100000 ; sin_tmp = 16'b0001000101000111 ; end 
  12'd140: begin cos_tmp = 16'b0011110110010010 ; sin_tmp = 16'b0001000101111000 ; end 
  12'd141: begin cos_tmp = 16'b0011110110010010 ; sin_tmp = 16'b0001000101111000 ; end 
  12'd142: begin cos_tmp = 16'b0011110110000100 ; sin_tmp = 16'b0001000110101010 ; end 
  12'd143: begin cos_tmp = 16'b0011110101110101 ; sin_tmp = 16'b0001000111011011 ; end 
  12'd144: begin cos_tmp = 16'b0011110101110101 ; sin_tmp = 16'b0001000111011011 ; end 
  12'd145: begin cos_tmp = 16'b0011110101100111 ; sin_tmp = 16'b0001001000001100 ; end 
  12'd146: begin cos_tmp = 16'b0011110101011000 ; sin_tmp = 16'b0001001000111110 ; end 
  12'd147: begin cos_tmp = 16'b0011110101011000 ; sin_tmp = 16'b0001001000111110 ; end 
  12'd148: begin cos_tmp = 16'b0011110101001010 ; sin_tmp = 16'b0001001001101111 ; end 
  12'd149: begin cos_tmp = 16'b0011110101001010 ; sin_tmp = 16'b0001001001101111 ; end 
  12'd150: begin cos_tmp = 16'b0011110100111011 ; sin_tmp = 16'b0001001010100000 ; end 
  12'd151: begin cos_tmp = 16'b0011110100101100 ; sin_tmp = 16'b0001001011010010 ; end 
  12'd152: begin cos_tmp = 16'b0011110100101100 ; sin_tmp = 16'b0001001011010010 ; end 
  12'd153: begin cos_tmp = 16'b0011110100011101 ; sin_tmp = 16'b0001001100000011 ; end 
  12'd154: begin cos_tmp = 16'b0011110100001101 ; sin_tmp = 16'b0001001100110100 ; end 
  12'd155: begin cos_tmp = 16'b0011110100001101 ; sin_tmp = 16'b0001001100110100 ; end 
  12'd156: begin cos_tmp = 16'b0011110011111110 ; sin_tmp = 16'b0001001101100101 ; end 
  12'd157: begin cos_tmp = 16'b0011110011111110 ; sin_tmp = 16'b0001001101100101 ; end 
  12'd158: begin cos_tmp = 16'b0011110011101110 ; sin_tmp = 16'b0001001110010110 ; end 
  12'd159: begin cos_tmp = 16'b0011110011011110 ; sin_tmp = 16'b0001001111000111 ; end 
  12'd160: begin cos_tmp = 16'b0011110011011110 ; sin_tmp = 16'b0001001111000111 ; end 
  12'd161: begin cos_tmp = 16'b0011110011001110 ; sin_tmp = 16'b0001001111111000 ; end 
  12'd162: begin cos_tmp = 16'b0011110010111110 ; sin_tmp = 16'b0001010000101001 ; end 
  12'd163: begin cos_tmp = 16'b0011110010111110 ; sin_tmp = 16'b0001010000101001 ; end 
  12'd164: begin cos_tmp = 16'b0011110010101110 ; sin_tmp = 16'b0001010001011010 ; end 
  12'd165: begin cos_tmp = 16'b0011110010101110 ; sin_tmp = 16'b0001010001011010 ; end 
  12'd166: begin cos_tmp = 16'b0011110010011101 ; sin_tmp = 16'b0001010010001010 ; end 
  12'd167: begin cos_tmp = 16'b0011110010001101 ; sin_tmp = 16'b0001010010111011 ; end 
  12'd168: begin cos_tmp = 16'b0011110010001101 ; sin_tmp = 16'b0001010010111011 ; end 
  12'd169: begin cos_tmp = 16'b0011110001111100 ; sin_tmp = 16'b0001010011101100 ; end 
  12'd170: begin cos_tmp = 16'b0011110001111100 ; sin_tmp = 16'b0001010011101100 ; end 
  12'd171: begin cos_tmp = 16'b0011110001101011 ; sin_tmp = 16'b0001010100011100 ; end 
  12'd172: begin cos_tmp = 16'b0011110001011010 ; sin_tmp = 16'b0001010101001101 ; end 
  12'd173: begin cos_tmp = 16'b0011110001011010 ; sin_tmp = 16'b0001010101001101 ; end 
  12'd174: begin cos_tmp = 16'b0011110001001001 ; sin_tmp = 16'b0001010101111101 ; end 
  12'd175: begin cos_tmp = 16'b0011110000110111 ; sin_tmp = 16'b0001010110101110 ; end 
  12'd176: begin cos_tmp = 16'b0011110000110111 ; sin_tmp = 16'b0001010110101110 ; end 
  12'd177: begin cos_tmp = 16'b0011110000100110 ; sin_tmp = 16'b0001010111011110 ; end 
  12'd178: begin cos_tmp = 16'b0011110000100110 ; sin_tmp = 16'b0001010111011110 ; end 
  12'd179: begin cos_tmp = 16'b0011110000010100 ; sin_tmp = 16'b0001011000001111 ; end 
  12'd180: begin cos_tmp = 16'b0011110000000010 ; sin_tmp = 16'b0001011000111111 ; end 
  12'd181: begin cos_tmp = 16'b0011110000000010 ; sin_tmp = 16'b0001011000111111 ; end 
  12'd182: begin cos_tmp = 16'b0011101111110000 ; sin_tmp = 16'b0001011001101111 ; end 
  12'd183: begin cos_tmp = 16'b0011101111011110 ; sin_tmp = 16'b0001011010011111 ; end 
  12'd184: begin cos_tmp = 16'b0011101111011110 ; sin_tmp = 16'b0001011010011111 ; end 
  12'd185: begin cos_tmp = 16'b0011101111001100 ; sin_tmp = 16'b0001011011001111 ; end 
  12'd186: begin cos_tmp = 16'b0011101111001100 ; sin_tmp = 16'b0001011011001111 ; end 
  12'd187: begin cos_tmp = 16'b0011101110111010 ; sin_tmp = 16'b0001011100000000 ; end 
  12'd188: begin cos_tmp = 16'b0011101110100111 ; sin_tmp = 16'b0001011100110000 ; end 
  12'd189: begin cos_tmp = 16'b0011101110100111 ; sin_tmp = 16'b0001011100110000 ; end 
  12'd190: begin cos_tmp = 16'b0011101110010100 ; sin_tmp = 16'b0001011101011111 ; end 
  12'd191: begin cos_tmp = 16'b0011101110000001 ; sin_tmp = 16'b0001011110001111 ; end 
  12'd192: begin cos_tmp = 16'b0011101110000001 ; sin_tmp = 16'b0001011110001111 ; end 
  12'd193: begin cos_tmp = 16'b0011101101101110 ; sin_tmp = 16'b0001011110111111 ; end 
  12'd194: begin cos_tmp = 16'b0011101101101110 ; sin_tmp = 16'b0001011110111111 ; end 
  12'd195: begin cos_tmp = 16'b0011101101011011 ; sin_tmp = 16'b0001011111101111 ; end 
  12'd196: begin cos_tmp = 16'b0011101101001000 ; sin_tmp = 16'b0001100000011111 ; end 
  12'd197: begin cos_tmp = 16'b0011101101001000 ; sin_tmp = 16'b0001100000011111 ; end 
  12'd198: begin cos_tmp = 16'b0011101100110100 ; sin_tmp = 16'b0001100001001110 ; end 
  12'd199: begin cos_tmp = 16'b0011101100100001 ; sin_tmp = 16'b0001100001111110 ; end 
  12'd200: begin cos_tmp = 16'b0011101100100001 ; sin_tmp = 16'b0001100001111110 ; end 
  12'd201: begin cos_tmp = 16'b0011101100001101 ; sin_tmp = 16'b0001100010101101 ; end 
  12'd202: begin cos_tmp = 16'b0011101100001101 ; sin_tmp = 16'b0001100010101101 ; end 
  12'd203: begin cos_tmp = 16'b0011101011111001 ; sin_tmp = 16'b0001100011011101 ; end 
  12'd204: begin cos_tmp = 16'b0011101011100101 ; sin_tmp = 16'b0001100100001100 ; end 
  12'd205: begin cos_tmp = 16'b0011101011100101 ; sin_tmp = 16'b0001100100001100 ; end 
  12'd206: begin cos_tmp = 16'b0011101011010001 ; sin_tmp = 16'b0001100100111100 ; end 
  12'd207: begin cos_tmp = 16'b0011101010111100 ; sin_tmp = 16'b0001100101101011 ; end 
  12'd208: begin cos_tmp = 16'b0011101010111100 ; sin_tmp = 16'b0001100101101011 ; end 
  12'd209: begin cos_tmp = 16'b0011101010101000 ; sin_tmp = 16'b0001100110011010 ; end 
  12'd210: begin cos_tmp = 16'b0011101010101000 ; sin_tmp = 16'b0001100110011010 ; end 
  12'd211: begin cos_tmp = 16'b0011101010010011 ; sin_tmp = 16'b0001100111001001 ; end 
  12'd212: begin cos_tmp = 16'b0011101001111110 ; sin_tmp = 16'b0001100111111000 ; end 
  12'd213: begin cos_tmp = 16'b0011101001111110 ; sin_tmp = 16'b0001100111111000 ; end 
  12'd214: begin cos_tmp = 16'b0011101001101010 ; sin_tmp = 16'b0001101000100111 ; end 
  12'd215: begin cos_tmp = 16'b0011101001101010 ; sin_tmp = 16'b0001101000100111 ; end 
  12'd216: begin cos_tmp = 16'b0011101001010100 ; sin_tmp = 16'b0001101001010110 ; end 
  12'd217: begin cos_tmp = 16'b0011101000111111 ; sin_tmp = 16'b0001101010000101 ; end 
  12'd218: begin cos_tmp = 16'b0011101000111111 ; sin_tmp = 16'b0001101010000101 ; end 
  12'd219: begin cos_tmp = 16'b0011101000101010 ; sin_tmp = 16'b0001101010110100 ; end 
  12'd220: begin cos_tmp = 16'b0011101000010100 ; sin_tmp = 16'b0001101011100011 ; end 
  12'd221: begin cos_tmp = 16'b0011101000010100 ; sin_tmp = 16'b0001101011100011 ; end 
  12'd222: begin cos_tmp = 16'b0011100111111111 ; sin_tmp = 16'b0001101100010001 ; end 
  12'd223: begin cos_tmp = 16'b0011100111111111 ; sin_tmp = 16'b0001101100010001 ; end 
  12'd224: begin cos_tmp = 16'b0011100111101001 ; sin_tmp = 16'b0001101101000000 ; end 
  12'd225: begin cos_tmp = 16'b0011100111010011 ; sin_tmp = 16'b0001101101101111 ; end 
  12'd226: begin cos_tmp = 16'b0011100111010011 ; sin_tmp = 16'b0001101101101111 ; end 
  12'd227: begin cos_tmp = 16'b0011100110111101 ; sin_tmp = 16'b0001101110011101 ; end 
  12'd228: begin cos_tmp = 16'b0011100110100110 ; sin_tmp = 16'b0001101111001011 ; end 
  12'd229: begin cos_tmp = 16'b0011100110100110 ; sin_tmp = 16'b0001101111001011 ; end 
  12'd230: begin cos_tmp = 16'b0011100110010000 ; sin_tmp = 16'b0001101111111010 ; end 
  12'd231: begin cos_tmp = 16'b0011100110010000 ; sin_tmp = 16'b0001101111111010 ; end 
  12'd232: begin cos_tmp = 16'b0011100101111001 ; sin_tmp = 16'b0001110000101000 ; end 
  12'd233: begin cos_tmp = 16'b0011100101100011 ; sin_tmp = 16'b0001110001010110 ; end 
  12'd234: begin cos_tmp = 16'b0011100101100011 ; sin_tmp = 16'b0001110001010110 ; end 
  12'd235: begin cos_tmp = 16'b0011100101001100 ; sin_tmp = 16'b0001110010000100 ; end 
  12'd236: begin cos_tmp = 16'b0011100100110101 ; sin_tmp = 16'b0001110010110010 ; end 
  12'd237: begin cos_tmp = 16'b0011100100110101 ; sin_tmp = 16'b0001110010110010 ; end 
  12'd238: begin cos_tmp = 16'b0011100100011110 ; sin_tmp = 16'b0001110011100000 ; end 
  12'd239: begin cos_tmp = 16'b0011100100011110 ; sin_tmp = 16'b0001110011100000 ; end 
  12'd240: begin cos_tmp = 16'b0011100100000110 ; sin_tmp = 16'b0001110100001110 ; end 
  12'd241: begin cos_tmp = 16'b0011100011101111 ; sin_tmp = 16'b0001110100111100 ; end 
  12'd242: begin cos_tmp = 16'b0011100011101111 ; sin_tmp = 16'b0001110100111100 ; end 
  12'd243: begin cos_tmp = 16'b0011100011010111 ; sin_tmp = 16'b0001110101101010 ; end 
  12'd244: begin cos_tmp = 16'b0011100011000000 ; sin_tmp = 16'b0001110110010111 ; end 
  12'd245: begin cos_tmp = 16'b0011100011000000 ; sin_tmp = 16'b0001110110010111 ; end 
  12'd246: begin cos_tmp = 16'b0011100010101000 ; sin_tmp = 16'b0001110111000101 ; end 
  12'd247: begin cos_tmp = 16'b0011100010101000 ; sin_tmp = 16'b0001110111000101 ; end 
  12'd248: begin cos_tmp = 16'b0011100010010000 ; sin_tmp = 16'b0001110111110011 ; end 
  12'd249: begin cos_tmp = 16'b0011100001110111 ; sin_tmp = 16'b0001111000100000 ; end 
  12'd250: begin cos_tmp = 16'b0011100001110111 ; sin_tmp = 16'b0001111000100000 ; end 
  12'd251: begin cos_tmp = 16'b0011100001011111 ; sin_tmp = 16'b0001111001001101 ; end 
  12'd252: begin cos_tmp = 16'b0011100001011111 ; sin_tmp = 16'b0001111001001101 ; end 
  12'd253: begin cos_tmp = 16'b0011100001000111 ; sin_tmp = 16'b0001111001111011 ; end 
  12'd254: begin cos_tmp = 16'b0011100000101110 ; sin_tmp = 16'b0001111010101000 ; end 
  12'd255: begin cos_tmp = 16'b0011100000101110 ; sin_tmp = 16'b0001111010101000 ; end 
  12'd256: begin cos_tmp = 16'b0011100000010101 ; sin_tmp = 16'b0001111011010101 ; end 
  12'd257: begin cos_tmp = 16'b0011011111111101 ; sin_tmp = 16'b0001111100000010 ; end 
  12'd258: begin cos_tmp = 16'b0011011111111101 ; sin_tmp = 16'b0001111100000010 ; end 
  12'd259: begin cos_tmp = 16'b0011011111100100 ; sin_tmp = 16'b0001111100101111 ; end 
  12'd260: begin cos_tmp = 16'b0011011111100100 ; sin_tmp = 16'b0001111100101111 ; end 
  12'd261: begin cos_tmp = 16'b0011011111001010 ; sin_tmp = 16'b0001111101011100 ; end 
  12'd262: begin cos_tmp = 16'b0011011110110001 ; sin_tmp = 16'b0001111110001001 ; end 
  12'd263: begin cos_tmp = 16'b0011011110110001 ; sin_tmp = 16'b0001111110001001 ; end 
  12'd264: begin cos_tmp = 16'b0011011110011000 ; sin_tmp = 16'b0001111110110110 ; end 
  12'd265: begin cos_tmp = 16'b0011011101111110 ; sin_tmp = 16'b0001111111100010 ; end 
  12'd266: begin cos_tmp = 16'b0011011101111110 ; sin_tmp = 16'b0001111111100010 ; end 
  12'd267: begin cos_tmp = 16'b0011011101100100 ; sin_tmp = 16'b0010000000001111 ; end 
  12'd268: begin cos_tmp = 16'b0011011101100100 ; sin_tmp = 16'b0010000000001111 ; end 
  12'd269: begin cos_tmp = 16'b0011011101001011 ; sin_tmp = 16'b0010000000111011 ; end 
  12'd270: begin cos_tmp = 16'b0011011100110001 ; sin_tmp = 16'b0010000001101000 ; end 
  12'd271: begin cos_tmp = 16'b0011011100110001 ; sin_tmp = 16'b0010000001101000 ; end 
  12'd272: begin cos_tmp = 16'b0011011100010110 ; sin_tmp = 16'b0010000010010100 ; end 
  12'd273: begin cos_tmp = 16'b0011011011111100 ; sin_tmp = 16'b0010000011000000 ; end 
  12'd274: begin cos_tmp = 16'b0011011011111100 ; sin_tmp = 16'b0010000011000000 ; end 
  12'd275: begin cos_tmp = 16'b0011011011100010 ; sin_tmp = 16'b0010000011101101 ; end 
  12'd276: begin cos_tmp = 16'b0011011011100010 ; sin_tmp = 16'b0010000011101101 ; end 
  12'd277: begin cos_tmp = 16'b0011011011000111 ; sin_tmp = 16'b0010000100011001 ; end 
  12'd278: begin cos_tmp = 16'b0011011010101100 ; sin_tmp = 16'b0010000101000101 ; end 
  12'd279: begin cos_tmp = 16'b0011011010101100 ; sin_tmp = 16'b0010000101000101 ; end 
  12'd280: begin cos_tmp = 16'b0011011010010010 ; sin_tmp = 16'b0010000101110001 ; end 
  12'd281: begin cos_tmp = 16'b0011011001110111 ; sin_tmp = 16'b0010000110011100 ; end 
  12'd282: begin cos_tmp = 16'b0011011001110111 ; sin_tmp = 16'b0010000110011100 ; end 
  12'd283: begin cos_tmp = 16'b0011011001011100 ; sin_tmp = 16'b0010000111001000 ; end 
  12'd284: begin cos_tmp = 16'b0011011001011100 ; sin_tmp = 16'b0010000111001000 ; end 
  12'd285: begin cos_tmp = 16'b0011011001000000 ; sin_tmp = 16'b0010000111110100 ; end 
  12'd286: begin cos_tmp = 16'b0011011000100101 ; sin_tmp = 16'b0010001000011111 ; end 
  12'd287: begin cos_tmp = 16'b0011011000100101 ; sin_tmp = 16'b0010001000011111 ; end 
  12'd288: begin cos_tmp = 16'b0011011000001001 ; sin_tmp = 16'b0010001001001011 ; end 
  12'd289: begin cos_tmp = 16'b0011011000001001 ; sin_tmp = 16'b0010001001001011 ; end 
  12'd290: begin cos_tmp = 16'b0011010111101110 ; sin_tmp = 16'b0010001001110110 ; end 
  12'd291: begin cos_tmp = 16'b0011010111010010 ; sin_tmp = 16'b0010001010100010 ; end 
  12'd292: begin cos_tmp = 16'b0011010111010010 ; sin_tmp = 16'b0010001010100010 ; end 
  12'd293: begin cos_tmp = 16'b0011010110110110 ; sin_tmp = 16'b0010001011001101 ; end 
  12'd294: begin cos_tmp = 16'b0011010110011010 ; sin_tmp = 16'b0010001011111000 ; end 
  12'd295: begin cos_tmp = 16'b0011010110011010 ; sin_tmp = 16'b0010001011111000 ; end 
  12'd296: begin cos_tmp = 16'b0011010101111110 ; sin_tmp = 16'b0010001100100011 ; end 
  12'd297: begin cos_tmp = 16'b0011010101111110 ; sin_tmp = 16'b0010001100100011 ; end 
  12'd298: begin cos_tmp = 16'b0011010101100010 ; sin_tmp = 16'b0010001101001110 ; end 
  12'd299: begin cos_tmp = 16'b0011010101000101 ; sin_tmp = 16'b0010001101111001 ; end 
  12'd300: begin cos_tmp = 16'b0011010101000101 ; sin_tmp = 16'b0010001101111001 ; end 
  12'd301: begin cos_tmp = 16'b0011010100101000 ; sin_tmp = 16'b0010001110100100 ; end 
  12'd302: begin cos_tmp = 16'b0011010100001100 ; sin_tmp = 16'b0010001111001111 ; end 
  12'd303: begin cos_tmp = 16'b0011010100001100 ; sin_tmp = 16'b0010001111001111 ; end 
  12'd304: begin cos_tmp = 16'b0011010011101111 ; sin_tmp = 16'b0010001111111001 ; end 
  12'd305: begin cos_tmp = 16'b0011010011101111 ; sin_tmp = 16'b0010001111111001 ; end 
  12'd306: begin cos_tmp = 16'b0011010011010010 ; sin_tmp = 16'b0010010000100100 ; end 
  12'd307: begin cos_tmp = 16'b0011010010110101 ; sin_tmp = 16'b0010010001001110 ; end 
  12'd308: begin cos_tmp = 16'b0011010010110101 ; sin_tmp = 16'b0010010001001110 ; end 
  12'd309: begin cos_tmp = 16'b0011010010010111 ; sin_tmp = 16'b0010010001111000 ; end 
  12'd310: begin cos_tmp = 16'b0011010001111010 ; sin_tmp = 16'b0010010010100011 ; end 
  12'd311: begin cos_tmp = 16'b0011010001111010 ; sin_tmp = 16'b0010010010100011 ; end 
  12'd312: begin cos_tmp = 16'b0011010001011101 ; sin_tmp = 16'b0010010011001101 ; end 
  12'd313: begin cos_tmp = 16'b0011010001011101 ; sin_tmp = 16'b0010010011001101 ; end 
  12'd314: begin cos_tmp = 16'b0011010000111111 ; sin_tmp = 16'b0010010011110111 ; end 
  12'd315: begin cos_tmp = 16'b0011010000100001 ; sin_tmp = 16'b0010010100100001 ; end 
  12'd316: begin cos_tmp = 16'b0011010000100001 ; sin_tmp = 16'b0010010100100001 ; end 
  12'd317: begin cos_tmp = 16'b0011010000000011 ; sin_tmp = 16'b0010010101001011 ; end 
  12'd318: begin cos_tmp = 16'b0011001111100101 ; sin_tmp = 16'b0010010101110101 ; end 
  12'd319: begin cos_tmp = 16'b0011001111100101 ; sin_tmp = 16'b0010010101110101 ; end 
  12'd320: begin cos_tmp = 16'b0011001111000111 ; sin_tmp = 16'b0010010110011110 ; end 
  12'd321: begin cos_tmp = 16'b0011001111000111 ; sin_tmp = 16'b0010010110011110 ; end 
  12'd322: begin cos_tmp = 16'b0011001110101001 ; sin_tmp = 16'b0010010111001000 ; end 
  12'd323: begin cos_tmp = 16'b0011001110001010 ; sin_tmp = 16'b0010010111110001 ; end 
  12'd324: begin cos_tmp = 16'b0011001110001010 ; sin_tmp = 16'b0010010111110001 ; end 
  12'd325: begin cos_tmp = 16'b0011001101101100 ; sin_tmp = 16'b0010011000011011 ; end 
  12'd326: begin cos_tmp = 16'b0011001101101100 ; sin_tmp = 16'b0010011000011011 ; end 
  12'd327: begin cos_tmp = 16'b0011001101001101 ; sin_tmp = 16'b0010011001000100 ; end 
  12'd328: begin cos_tmp = 16'b0011001100101110 ; sin_tmp = 16'b0010011001101101 ; end 
  12'd329: begin cos_tmp = 16'b0011001100101110 ; sin_tmp = 16'b0010011001101101 ; end 
  12'd330: begin cos_tmp = 16'b0011001100001111 ; sin_tmp = 16'b0010011010010110 ; end 
  12'd331: begin cos_tmp = 16'b0011001011110000 ; sin_tmp = 16'b0010011010111111 ; end 
  12'd332: begin cos_tmp = 16'b0011001011110000 ; sin_tmp = 16'b0010011010111111 ; end 
  12'd333: begin cos_tmp = 16'b0011001011010001 ; sin_tmp = 16'b0010011011101000 ; end 
  12'd334: begin cos_tmp = 16'b0011001011010001 ; sin_tmp = 16'b0010011011101000 ; end 
  12'd335: begin cos_tmp = 16'b0011001010110001 ; sin_tmp = 16'b0010011100010001 ; end 
  12'd336: begin cos_tmp = 16'b0011001010010010 ; sin_tmp = 16'b0010011100111010 ; end 
  12'd337: begin cos_tmp = 16'b0011001010010010 ; sin_tmp = 16'b0010011100111010 ; end 
  12'd338: begin cos_tmp = 16'b0011001001110010 ; sin_tmp = 16'b0010011101100010 ; end 
  12'd339: begin cos_tmp = 16'b0011001001010011 ; sin_tmp = 16'b0010011110001011 ; end 
  12'd340: begin cos_tmp = 16'b0011001001010011 ; sin_tmp = 16'b0010011110001011 ; end 
  12'd341: begin cos_tmp = 16'b0011001000110011 ; sin_tmp = 16'b0010011110110011 ; end 
  12'd342: begin cos_tmp = 16'b0011001000110011 ; sin_tmp = 16'b0010011110110011 ; end 
  12'd343: begin cos_tmp = 16'b0011001000010011 ; sin_tmp = 16'b0010011111011100 ; end 
  12'd344: begin cos_tmp = 16'b0011000111110011 ; sin_tmp = 16'b0010100000000100 ; end 
  12'd345: begin cos_tmp = 16'b0011000111110011 ; sin_tmp = 16'b0010100000000100 ; end 
  12'd346: begin cos_tmp = 16'b0011000111010010 ; sin_tmp = 16'b0010100000101100 ; end 
  12'd347: begin cos_tmp = 16'b0011000110110010 ; sin_tmp = 16'b0010100001010100 ; end 
  12'd348: begin cos_tmp = 16'b0011000110110010 ; sin_tmp = 16'b0010100001010100 ; end 
  12'd349: begin cos_tmp = 16'b0011000110010001 ; sin_tmp = 16'b0010100001111100 ; end 
  12'd350: begin cos_tmp = 16'b0011000110010001 ; sin_tmp = 16'b0010100001111100 ; end 
  12'd351: begin cos_tmp = 16'b0011000101110001 ; sin_tmp = 16'b0010100010100100 ; end 
  12'd352: begin cos_tmp = 16'b0011000101010000 ; sin_tmp = 16'b0010100011001100 ; end 
  12'd353: begin cos_tmp = 16'b0011000101010000 ; sin_tmp = 16'b0010100011001100 ; end 
  12'd354: begin cos_tmp = 16'b0011000100101111 ; sin_tmp = 16'b0010100011110011 ; end 
  12'd355: begin cos_tmp = 16'b0011000100001110 ; sin_tmp = 16'b0010100100011011 ; end 
  12'd356: begin cos_tmp = 16'b0011000100001110 ; sin_tmp = 16'b0010100100011011 ; end 
  12'd357: begin cos_tmp = 16'b0011000011101101 ; sin_tmp = 16'b0010100101000010 ; end 
  12'd358: begin cos_tmp = 16'b0011000011101101 ; sin_tmp = 16'b0010100101000010 ; end 
  12'd359: begin cos_tmp = 16'b0011000011001100 ; sin_tmp = 16'b0010100101101001 ; end 
  12'd360: begin cos_tmp = 16'b0011000010101010 ; sin_tmp = 16'b0010100110010001 ; end 
  12'd361: begin cos_tmp = 16'b0011000010101010 ; sin_tmp = 16'b0010100110010001 ; end 
  12'd362: begin cos_tmp = 16'b0011000010001001 ; sin_tmp = 16'b0010100110111000 ; end 
  12'd363: begin cos_tmp = 16'b0011000010001001 ; sin_tmp = 16'b0010100110111000 ; end 
  12'd364: begin cos_tmp = 16'b0011000001100111 ; sin_tmp = 16'b0010100111011111 ; end 
  12'd365: begin cos_tmp = 16'b0011000001000110 ; sin_tmp = 16'b0010101000000110 ; end 
  12'd366: begin cos_tmp = 16'b0011000001000110 ; sin_tmp = 16'b0010101000000110 ; end 
  12'd367: begin cos_tmp = 16'b0011000000100100 ; sin_tmp = 16'b0010101000101100 ; end 
  12'd368: begin cos_tmp = 16'b0011000000000010 ; sin_tmp = 16'b0010101001010011 ; end 
  12'd369: begin cos_tmp = 16'b0011000000000010 ; sin_tmp = 16'b0010101001010011 ; end 
  12'd370: begin cos_tmp = 16'b0010111111100000 ; sin_tmp = 16'b0010101001111001 ; end 
  12'd371: begin cos_tmp = 16'b0010111111100000 ; sin_tmp = 16'b0010101001111001 ; end 
  12'd372: begin cos_tmp = 16'b0010111110111101 ; sin_tmp = 16'b0010101010100000 ; end 
  12'd373: begin cos_tmp = 16'b0010111110011011 ; sin_tmp = 16'b0010101011000110 ; end 
  12'd374: begin cos_tmp = 16'b0010111110011011 ; sin_tmp = 16'b0010101011000110 ; end 
  12'd375: begin cos_tmp = 16'b0010111101111001 ; sin_tmp = 16'b0010101011101101 ; end 
  12'd376: begin cos_tmp = 16'b0010111101010110 ; sin_tmp = 16'b0010101100010011 ; end 
  12'd377: begin cos_tmp = 16'b0010111101010110 ; sin_tmp = 16'b0010101100010011 ; end 
  12'd378: begin cos_tmp = 16'b0010111100110011 ; sin_tmp = 16'b0010101100111001 ; end 
  12'd379: begin cos_tmp = 16'b0010111100110011 ; sin_tmp = 16'b0010101100111001 ; end 
  12'd380: begin cos_tmp = 16'b0010111100010001 ; sin_tmp = 16'b0010101101011111 ; end 
  12'd381: begin cos_tmp = 16'b0010111011101110 ; sin_tmp = 16'b0010101110000100 ; end 
  12'd382: begin cos_tmp = 16'b0010111011101110 ; sin_tmp = 16'b0010101110000100 ; end 
  12'd383: begin cos_tmp = 16'b0010111011001011 ; sin_tmp = 16'b0010101110101010 ; end 
  12'd384: begin cos_tmp = 16'b0010111010100111 ; sin_tmp = 16'b0010101111010000 ; end 
  12'd385: begin cos_tmp = 16'b0010111010100111 ; sin_tmp = 16'b0010101111010000 ; end 
  12'd386: begin cos_tmp = 16'b0010111010000100 ; sin_tmp = 16'b0010101111110101 ; end 
  12'd387: begin cos_tmp = 16'b0010111010000100 ; sin_tmp = 16'b0010101111110101 ; end 
  12'd388: begin cos_tmp = 16'b0010111001100001 ; sin_tmp = 16'b0010110000011010 ; end 
  12'd389: begin cos_tmp = 16'b0010111000111101 ; sin_tmp = 16'b0010110001000000 ; end 
  12'd390: begin cos_tmp = 16'b0010111000111101 ; sin_tmp = 16'b0010110001000000 ; end 
  12'd391: begin cos_tmp = 16'b0010111000011010 ; sin_tmp = 16'b0010110001100101 ; end 
  12'd392: begin cos_tmp = 16'b0010110111110110 ; sin_tmp = 16'b0010110010001010 ; end 
  12'd393: begin cos_tmp = 16'b0010110111110110 ; sin_tmp = 16'b0010110010001010 ; end 
  12'd394: begin cos_tmp = 16'b0010110111010010 ; sin_tmp = 16'b0010110010101111 ; end 
  12'd395: begin cos_tmp = 16'b0010110111010010 ; sin_tmp = 16'b0010110010101111 ; end 
  12'd396: begin cos_tmp = 16'b0010110110101110 ; sin_tmp = 16'b0010110011010100 ; end 
  12'd397: begin cos_tmp = 16'b0010110110001010 ; sin_tmp = 16'b0010110011111000 ; end 
  12'd398: begin cos_tmp = 16'b0010110110001010 ; sin_tmp = 16'b0010110011111000 ; end 
  12'd399: begin cos_tmp = 16'b0010110101100110 ; sin_tmp = 16'b0010110100011101 ; end 
  12'd400: begin cos_tmp = 16'b0010110101100110 ; sin_tmp = 16'b0010110100011101 ; end 
  12'd401: begin cos_tmp = 16'b0010110101000001 ; sin_tmp = 16'b0010110101000001 ; end 
  12'd402: begin cos_tmp = 16'b0010110100011101 ; sin_tmp = 16'b0010110101100110 ; end 
  12'd403: begin cos_tmp = 16'b0010110100011101 ; sin_tmp = 16'b0010110101100110 ; end 
  12'd404: begin cos_tmp = 16'b0010110011111000 ; sin_tmp = 16'b0010110110001010 ; end 
  12'd405: begin cos_tmp = 16'b0010110011010100 ; sin_tmp = 16'b0010110110101110 ; end 
  12'd406: begin cos_tmp = 16'b0010110011010100 ; sin_tmp = 16'b0010110110101110 ; end 
  12'd407: begin cos_tmp = 16'b0010110010101111 ; sin_tmp = 16'b0010110111010010 ; end 
  12'd408: begin cos_tmp = 16'b0010110010101111 ; sin_tmp = 16'b0010110111010010 ; end 
  12'd409: begin cos_tmp = 16'b0010110010001010 ; sin_tmp = 16'b0010110111110110 ; end 
  12'd410: begin cos_tmp = 16'b0010110001100101 ; sin_tmp = 16'b0010111000011010 ; end 
  12'd411: begin cos_tmp = 16'b0010110001100101 ; sin_tmp = 16'b0010111000011010 ; end 
  12'd412: begin cos_tmp = 16'b0010110001000000 ; sin_tmp = 16'b0010111000111101 ; end 
  12'd413: begin cos_tmp = 16'b0010110000011010 ; sin_tmp = 16'b0010111001100001 ; end 
  12'd414: begin cos_tmp = 16'b0010110000011010 ; sin_tmp = 16'b0010111001100001 ; end 
  12'd415: begin cos_tmp = 16'b0010101111110101 ; sin_tmp = 16'b0010111010000100 ; end 
  12'd416: begin cos_tmp = 16'b0010101111110101 ; sin_tmp = 16'b0010111010000100 ; end 
  12'd417: begin cos_tmp = 16'b0010101111010000 ; sin_tmp = 16'b0010111010100111 ; end 
  12'd418: begin cos_tmp = 16'b0010101110101010 ; sin_tmp = 16'b0010111011001011 ; end 
  12'd419: begin cos_tmp = 16'b0010101110101010 ; sin_tmp = 16'b0010111011001011 ; end 
  12'd420: begin cos_tmp = 16'b0010101110000100 ; sin_tmp = 16'b0010111011101110 ; end 
  12'd421: begin cos_tmp = 16'b0010101101011111 ; sin_tmp = 16'b0010111100010001 ; end 
  12'd422: begin cos_tmp = 16'b0010101101011111 ; sin_tmp = 16'b0010111100010001 ; end 
  12'd423: begin cos_tmp = 16'b0010101100111001 ; sin_tmp = 16'b0010111100110011 ; end 
  12'd424: begin cos_tmp = 16'b0010101100111001 ; sin_tmp = 16'b0010111100110011 ; end 
  12'd425: begin cos_tmp = 16'b0010101100010011 ; sin_tmp = 16'b0010111101010110 ; end 
  12'd426: begin cos_tmp = 16'b0010101011101101 ; sin_tmp = 16'b0010111101111001 ; end 
  12'd427: begin cos_tmp = 16'b0010101011101101 ; sin_tmp = 16'b0010111101111001 ; end 
  12'd428: begin cos_tmp = 16'b0010101011000110 ; sin_tmp = 16'b0010111110011011 ; end 
  12'd429: begin cos_tmp = 16'b0010101010100000 ; sin_tmp = 16'b0010111110111101 ; end 
  12'd430: begin cos_tmp = 16'b0010101010100000 ; sin_tmp = 16'b0010111110111101 ; end 
  12'd431: begin cos_tmp = 16'b0010101001111001 ; sin_tmp = 16'b0010111111100000 ; end 
  12'd432: begin cos_tmp = 16'b0010101001111001 ; sin_tmp = 16'b0010111111100000 ; end 
  12'd433: begin cos_tmp = 16'b0010101001010011 ; sin_tmp = 16'b0011000000000010 ; end 
  12'd434: begin cos_tmp = 16'b0010101000101100 ; sin_tmp = 16'b0011000000100100 ; end 
  12'd435: begin cos_tmp = 16'b0010101000101100 ; sin_tmp = 16'b0011000000100100 ; end 
  12'd436: begin cos_tmp = 16'b0010101000000110 ; sin_tmp = 16'b0011000001000110 ; end 
  12'd437: begin cos_tmp = 16'b0010101000000110 ; sin_tmp = 16'b0011000001000110 ; end 
  12'd438: begin cos_tmp = 16'b0010100111011111 ; sin_tmp = 16'b0011000001100111 ; end 
  12'd439: begin cos_tmp = 16'b0010100110111000 ; sin_tmp = 16'b0011000010001001 ; end 
  12'd440: begin cos_tmp = 16'b0010100110111000 ; sin_tmp = 16'b0011000010001001 ; end 
  12'd441: begin cos_tmp = 16'b0010100110010001 ; sin_tmp = 16'b0011000010101010 ; end 
  12'd442: begin cos_tmp = 16'b0010100101101001 ; sin_tmp = 16'b0011000011001100 ; end 
  12'd443: begin cos_tmp = 16'b0010100101101001 ; sin_tmp = 16'b0011000011001100 ; end 
  12'd444: begin cos_tmp = 16'b0010100101000010 ; sin_tmp = 16'b0011000011101101 ; end 
  12'd445: begin cos_tmp = 16'b0010100101000010 ; sin_tmp = 16'b0011000011101101 ; end 
  12'd446: begin cos_tmp = 16'b0010100100011011 ; sin_tmp = 16'b0011000100001110 ; end 
  12'd447: begin cos_tmp = 16'b0010100011110011 ; sin_tmp = 16'b0011000100101111 ; end 
  12'd448: begin cos_tmp = 16'b0010100011110011 ; sin_tmp = 16'b0011000100101111 ; end 
  12'd449: begin cos_tmp = 16'b0010100011001100 ; sin_tmp = 16'b0011000101010000 ; end 
  12'd450: begin cos_tmp = 16'b0010100010100100 ; sin_tmp = 16'b0011000101110001 ; end 
  12'd451: begin cos_tmp = 16'b0010100010100100 ; sin_tmp = 16'b0011000101110001 ; end 
  12'd452: begin cos_tmp = 16'b0010100001111100 ; sin_tmp = 16'b0011000110010001 ; end 
  12'd453: begin cos_tmp = 16'b0010100001111100 ; sin_tmp = 16'b0011000110010001 ; end 
  12'd454: begin cos_tmp = 16'b0010100001010100 ; sin_tmp = 16'b0011000110110010 ; end 
  12'd455: begin cos_tmp = 16'b0010100000101100 ; sin_tmp = 16'b0011000111010010 ; end 
  12'd456: begin cos_tmp = 16'b0010100000101100 ; sin_tmp = 16'b0011000111010010 ; end 
  12'd457: begin cos_tmp = 16'b0010100000000100 ; sin_tmp = 16'b0011000111110011 ; end 
  12'd458: begin cos_tmp = 16'b0010011111011100 ; sin_tmp = 16'b0011001000010011 ; end 
  12'd459: begin cos_tmp = 16'b0010011111011100 ; sin_tmp = 16'b0011001000010011 ; end 
  12'd460: begin cos_tmp = 16'b0010011110110011 ; sin_tmp = 16'b0011001000110011 ; end 
  12'd461: begin cos_tmp = 16'b0010011110110011 ; sin_tmp = 16'b0011001000110011 ; end 
  12'd462: begin cos_tmp = 16'b0010011110001011 ; sin_tmp = 16'b0011001001010011 ; end 
  12'd463: begin cos_tmp = 16'b0010011101100010 ; sin_tmp = 16'b0011001001110010 ; end 
  12'd464: begin cos_tmp = 16'b0010011101100010 ; sin_tmp = 16'b0011001001110010 ; end 
  12'd465: begin cos_tmp = 16'b0010011100111010 ; sin_tmp = 16'b0011001010010010 ; end 
  12'd466: begin cos_tmp = 16'b0010011100010001 ; sin_tmp = 16'b0011001010110001 ; end 
  12'd467: begin cos_tmp = 16'b0010011100010001 ; sin_tmp = 16'b0011001010110001 ; end 
  12'd468: begin cos_tmp = 16'b0010011011101000 ; sin_tmp = 16'b0011001011010001 ; end 
  12'd469: begin cos_tmp = 16'b0010011011101000 ; sin_tmp = 16'b0011001011010001 ; end 
  12'd470: begin cos_tmp = 16'b0010011010111111 ; sin_tmp = 16'b0011001011110000 ; end 
  12'd471: begin cos_tmp = 16'b0010011010010110 ; sin_tmp = 16'b0011001100001111 ; end 
  12'd472: begin cos_tmp = 16'b0010011010010110 ; sin_tmp = 16'b0011001100001111 ; end 
  12'd473: begin cos_tmp = 16'b0010011001101101 ; sin_tmp = 16'b0011001100101110 ; end 
  12'd474: begin cos_tmp = 16'b0010011001101101 ; sin_tmp = 16'b0011001100101110 ; end 
  12'd475: begin cos_tmp = 16'b0010011001000100 ; sin_tmp = 16'b0011001101001101 ; end 
  12'd476: begin cos_tmp = 16'b0010011000011011 ; sin_tmp = 16'b0011001101101100 ; end 
  12'd477: begin cos_tmp = 16'b0010011000011011 ; sin_tmp = 16'b0011001101101100 ; end 
  12'd478: begin cos_tmp = 16'b0010010111110001 ; sin_tmp = 16'b0011001110001010 ; end 
  12'd479: begin cos_tmp = 16'b0010010111001000 ; sin_tmp = 16'b0011001110101001 ; end 
  12'd480: begin cos_tmp = 16'b0010010111001000 ; sin_tmp = 16'b0011001110101001 ; end 
  12'd481: begin cos_tmp = 16'b0010010110011110 ; sin_tmp = 16'b0011001111000111 ; end 
  12'd482: begin cos_tmp = 16'b0010010110011110 ; sin_tmp = 16'b0011001111000111 ; end 
  12'd483: begin cos_tmp = 16'b0010010101110101 ; sin_tmp = 16'b0011001111100101 ; end 
  12'd484: begin cos_tmp = 16'b0010010101001011 ; sin_tmp = 16'b0011010000000011 ; end 
  12'd485: begin cos_tmp = 16'b0010010101001011 ; sin_tmp = 16'b0011010000000011 ; end 
  12'd486: begin cos_tmp = 16'b0010010100100001 ; sin_tmp = 16'b0011010000100001 ; end 
  12'd487: begin cos_tmp = 16'b0010010011110111 ; sin_tmp = 16'b0011010000111111 ; end 
  12'd488: begin cos_tmp = 16'b0010010011110111 ; sin_tmp = 16'b0011010000111111 ; end 
  12'd489: begin cos_tmp = 16'b0010010011001101 ; sin_tmp = 16'b0011010001011101 ; end 
  12'd490: begin cos_tmp = 16'b0010010011001101 ; sin_tmp = 16'b0011010001011101 ; end 
  12'd491: begin cos_tmp = 16'b0010010010100011 ; sin_tmp = 16'b0011010001111010 ; end 
  12'd492: begin cos_tmp = 16'b0010010001111000 ; sin_tmp = 16'b0011010010010111 ; end 
  12'd493: begin cos_tmp = 16'b0010010001111000 ; sin_tmp = 16'b0011010010010111 ; end 
  12'd494: begin cos_tmp = 16'b0010010001001110 ; sin_tmp = 16'b0011010010110101 ; end 
  12'd495: begin cos_tmp = 16'b0010010000100100 ; sin_tmp = 16'b0011010011010010 ; end 
  12'd496: begin cos_tmp = 16'b0010010000100100 ; sin_tmp = 16'b0011010011010010 ; end 
  12'd497: begin cos_tmp = 16'b0010001111111001 ; sin_tmp = 16'b0011010011101111 ; end 
  12'd498: begin cos_tmp = 16'b0010001111111001 ; sin_tmp = 16'b0011010011101111 ; end 
  12'd499: begin cos_tmp = 16'b0010001111001111 ; sin_tmp = 16'b0011010100001100 ; end 
  12'd500: begin cos_tmp = 16'b0010001110100100 ; sin_tmp = 16'b0011010100101000 ; end 
  12'd501: begin cos_tmp = 16'b0010001110100100 ; sin_tmp = 16'b0011010100101000 ; end 
  12'd502: begin cos_tmp = 16'b0010001101111001 ; sin_tmp = 16'b0011010101000101 ; end 
  12'd503: begin cos_tmp = 16'b0010001101001110 ; sin_tmp = 16'b0011010101100010 ; end 
  12'd504: begin cos_tmp = 16'b0010001101001110 ; sin_tmp = 16'b0011010101100010 ; end 
  12'd505: begin cos_tmp = 16'b0010001100100011 ; sin_tmp = 16'b0011010101111110 ; end 
  12'd506: begin cos_tmp = 16'b0010001100100011 ; sin_tmp = 16'b0011010101111110 ; end 
  12'd507: begin cos_tmp = 16'b0010001011111000 ; sin_tmp = 16'b0011010110011010 ; end 
  12'd508: begin cos_tmp = 16'b0010001011001101 ; sin_tmp = 16'b0011010110110110 ; end 
  12'd509: begin cos_tmp = 16'b0010001011001101 ; sin_tmp = 16'b0011010110110110 ; end 
  12'd510: begin cos_tmp = 16'b0010001010100010 ; sin_tmp = 16'b0011010111010010 ; end 
  12'd511: begin cos_tmp = 16'b0010001010100010 ; sin_tmp = 16'b0011010111010010 ; end 
  12'd512: begin cos_tmp = 16'b0010001001110110 ; sin_tmp = 16'b0011010111101110 ; end 
  12'd513: begin cos_tmp = 16'b0010001001001011 ; sin_tmp = 16'b0011011000001001 ; end 
  12'd514: begin cos_tmp = 16'b0010001001001011 ; sin_tmp = 16'b0011011000001001 ; end 
  12'd515: begin cos_tmp = 16'b0010001000011111 ; sin_tmp = 16'b0011011000100101 ; end 
  12'd516: begin cos_tmp = 16'b0010000111110100 ; sin_tmp = 16'b0011011001000000 ; end 
  12'd517: begin cos_tmp = 16'b0010000111110100 ; sin_tmp = 16'b0011011001000000 ; end 
  12'd518: begin cos_tmp = 16'b0010000111001000 ; sin_tmp = 16'b0011011001011100 ; end 
  12'd519: begin cos_tmp = 16'b0010000111001000 ; sin_tmp = 16'b0011011001011100 ; end 
  12'd520: begin cos_tmp = 16'b0010000110011100 ; sin_tmp = 16'b0011011001110111 ; end 
  12'd521: begin cos_tmp = 16'b0010000101110001 ; sin_tmp = 16'b0011011010010010 ; end 
  12'd522: begin cos_tmp = 16'b0010000101110001 ; sin_tmp = 16'b0011011010010010 ; end 
  12'd523: begin cos_tmp = 16'b0010000101000101 ; sin_tmp = 16'b0011011010101100 ; end 
  12'd524: begin cos_tmp = 16'b0010000100011001 ; sin_tmp = 16'b0011011011000111 ; end 
  12'd525: begin cos_tmp = 16'b0010000100011001 ; sin_tmp = 16'b0011011011000111 ; end 
  12'd526: begin cos_tmp = 16'b0010000011101101 ; sin_tmp = 16'b0011011011100010 ; end 
  12'd527: begin cos_tmp = 16'b0010000011101101 ; sin_tmp = 16'b0011011011100010 ; end 
  12'd528: begin cos_tmp = 16'b0010000011000000 ; sin_tmp = 16'b0011011011111100 ; end 
  12'd529: begin cos_tmp = 16'b0010000010010100 ; sin_tmp = 16'b0011011100010110 ; end 
  12'd530: begin cos_tmp = 16'b0010000010010100 ; sin_tmp = 16'b0011011100010110 ; end 
  12'd531: begin cos_tmp = 16'b0010000001101000 ; sin_tmp = 16'b0011011100110001 ; end 
  12'd532: begin cos_tmp = 16'b0010000000111011 ; sin_tmp = 16'b0011011101001011 ; end 
  12'd533: begin cos_tmp = 16'b0010000000111011 ; sin_tmp = 16'b0011011101001011 ; end 
  12'd534: begin cos_tmp = 16'b0010000000001111 ; sin_tmp = 16'b0011011101100100 ; end 
  12'd535: begin cos_tmp = 16'b0010000000001111 ; sin_tmp = 16'b0011011101100100 ; end 
  12'd536: begin cos_tmp = 16'b0001111111100010 ; sin_tmp = 16'b0011011101111110 ; end 
  12'd537: begin cos_tmp = 16'b0001111110110110 ; sin_tmp = 16'b0011011110011000 ; end 
  12'd538: begin cos_tmp = 16'b0001111110110110 ; sin_tmp = 16'b0011011110011000 ; end 
  12'd539: begin cos_tmp = 16'b0001111110001001 ; sin_tmp = 16'b0011011110110001 ; end 
  12'd540: begin cos_tmp = 16'b0001111101011100 ; sin_tmp = 16'b0011011111001010 ; end 
  12'd541: begin cos_tmp = 16'b0001111101011100 ; sin_tmp = 16'b0011011111001010 ; end 
  12'd542: begin cos_tmp = 16'b0001111100101111 ; sin_tmp = 16'b0011011111100100 ; end 
  12'd543: begin cos_tmp = 16'b0001111100101111 ; sin_tmp = 16'b0011011111100100 ; end 
  12'd544: begin cos_tmp = 16'b0001111100000010 ; sin_tmp = 16'b0011011111111101 ; end 
  12'd545: begin cos_tmp = 16'b0001111011010101 ; sin_tmp = 16'b0011100000010101 ; end 
  12'd546: begin cos_tmp = 16'b0001111011010101 ; sin_tmp = 16'b0011100000010101 ; end 
  12'd547: begin cos_tmp = 16'b0001111010101000 ; sin_tmp = 16'b0011100000101110 ; end 
  12'd548: begin cos_tmp = 16'b0001111001111011 ; sin_tmp = 16'b0011100001000111 ; end 
  12'd549: begin cos_tmp = 16'b0001111001111011 ; sin_tmp = 16'b0011100001000111 ; end 
  12'd550: begin cos_tmp = 16'b0001111001001101 ; sin_tmp = 16'b0011100001011111 ; end 
  12'd551: begin cos_tmp = 16'b0001111001001101 ; sin_tmp = 16'b0011100001011111 ; end 
  12'd552: begin cos_tmp = 16'b0001111000100000 ; sin_tmp = 16'b0011100001110111 ; end 
  12'd553: begin cos_tmp = 16'b0001110111110011 ; sin_tmp = 16'b0011100010010000 ; end 
  12'd554: begin cos_tmp = 16'b0001110111110011 ; sin_tmp = 16'b0011100010010000 ; end 
  12'd555: begin cos_tmp = 16'b0001110111000101 ; sin_tmp = 16'b0011100010101000 ; end 
  12'd556: begin cos_tmp = 16'b0001110111000101 ; sin_tmp = 16'b0011100010101000 ; end 
  12'd557: begin cos_tmp = 16'b0001110110010111 ; sin_tmp = 16'b0011100011000000 ; end 
  12'd558: begin cos_tmp = 16'b0001110101101010 ; sin_tmp = 16'b0011100011010111 ; end 
  12'd559: begin cos_tmp = 16'b0001110101101010 ; sin_tmp = 16'b0011100011010111 ; end 
  12'd560: begin cos_tmp = 16'b0001110100111100 ; sin_tmp = 16'b0011100011101111 ; end 
  12'd561: begin cos_tmp = 16'b0001110100001110 ; sin_tmp = 16'b0011100100000110 ; end 
  12'd562: begin cos_tmp = 16'b0001110100001110 ; sin_tmp = 16'b0011100100000110 ; end 
  12'd563: begin cos_tmp = 16'b0001110011100000 ; sin_tmp = 16'b0011100100011110 ; end 
  12'd564: begin cos_tmp = 16'b0001110011100000 ; sin_tmp = 16'b0011100100011110 ; end 
  12'd565: begin cos_tmp = 16'b0001110010110010 ; sin_tmp = 16'b0011100100110101 ; end 
  12'd566: begin cos_tmp = 16'b0001110010000100 ; sin_tmp = 16'b0011100101001100 ; end 
  12'd567: begin cos_tmp = 16'b0001110010000100 ; sin_tmp = 16'b0011100101001100 ; end 
  12'd568: begin cos_tmp = 16'b0001110001010110 ; sin_tmp = 16'b0011100101100011 ; end 
  12'd569: begin cos_tmp = 16'b0001110000101000 ; sin_tmp = 16'b0011100101111001 ; end 
  12'd570: begin cos_tmp = 16'b0001110000101000 ; sin_tmp = 16'b0011100101111001 ; end 
  12'd571: begin cos_tmp = 16'b0001101111111010 ; sin_tmp = 16'b0011100110010000 ; end 
  12'd572: begin cos_tmp = 16'b0001101111111010 ; sin_tmp = 16'b0011100110010000 ; end 
  12'd573: begin cos_tmp = 16'b0001101111001011 ; sin_tmp = 16'b0011100110100110 ; end 
  12'd574: begin cos_tmp = 16'b0001101110011101 ; sin_tmp = 16'b0011100110111101 ; end 
  12'd575: begin cos_tmp = 16'b0001101110011101 ; sin_tmp = 16'b0011100110111101 ; end 
  12'd576: begin cos_tmp = 16'b0001101101101111 ; sin_tmp = 16'b0011100111010011 ; end 
  12'd577: begin cos_tmp = 16'b0001101101000000 ; sin_tmp = 16'b0011100111101001 ; end 
  12'd578: begin cos_tmp = 16'b0001101101000000 ; sin_tmp = 16'b0011100111101001 ; end 
  12'd579: begin cos_tmp = 16'b0001101100010001 ; sin_tmp = 16'b0011100111111111 ; end 
  12'd580: begin cos_tmp = 16'b0001101100010001 ; sin_tmp = 16'b0011100111111111 ; end 
  12'd581: begin cos_tmp = 16'b0001101011100011 ; sin_tmp = 16'b0011101000010100 ; end 
  12'd582: begin cos_tmp = 16'b0001101010110100 ; sin_tmp = 16'b0011101000101010 ; end 
  12'd583: begin cos_tmp = 16'b0001101010110100 ; sin_tmp = 16'b0011101000101010 ; end 
  12'd584: begin cos_tmp = 16'b0001101010000101 ; sin_tmp = 16'b0011101000111111 ; end 
  12'd585: begin cos_tmp = 16'b0001101001010110 ; sin_tmp = 16'b0011101001010100 ; end 
  12'd586: begin cos_tmp = 16'b0001101001010110 ; sin_tmp = 16'b0011101001010100 ; end 
  12'd587: begin cos_tmp = 16'b0001101000100111 ; sin_tmp = 16'b0011101001101010 ; end 
  12'd588: begin cos_tmp = 16'b0001101000100111 ; sin_tmp = 16'b0011101001101010 ; end 
  12'd589: begin cos_tmp = 16'b0001100111111000 ; sin_tmp = 16'b0011101001111110 ; end 
  12'd590: begin cos_tmp = 16'b0001100111001001 ; sin_tmp = 16'b0011101010010011 ; end 
  12'd591: begin cos_tmp = 16'b0001100111001001 ; sin_tmp = 16'b0011101010010011 ; end 
  12'd592: begin cos_tmp = 16'b0001100110011010 ; sin_tmp = 16'b0011101010101000 ; end 
  12'd593: begin cos_tmp = 16'b0001100110011010 ; sin_tmp = 16'b0011101010101000 ; end 
  12'd594: begin cos_tmp = 16'b0001100101101011 ; sin_tmp = 16'b0011101010111100 ; end 
  12'd595: begin cos_tmp = 16'b0001100100111100 ; sin_tmp = 16'b0011101011010001 ; end 
  12'd596: begin cos_tmp = 16'b0001100100111100 ; sin_tmp = 16'b0011101011010001 ; end 
  12'd597: begin cos_tmp = 16'b0001100100001100 ; sin_tmp = 16'b0011101011100101 ; end 
  12'd598: begin cos_tmp = 16'b0001100011011101 ; sin_tmp = 16'b0011101011111001 ; end 
  12'd599: begin cos_tmp = 16'b0001100011011101 ; sin_tmp = 16'b0011101011111001 ; end 
  12'd600: begin cos_tmp = 16'b0001100010101101 ; sin_tmp = 16'b0011101100001101 ; end 
  12'd601: begin cos_tmp = 16'b0001100010101101 ; sin_tmp = 16'b0011101100001101 ; end 
  12'd602: begin cos_tmp = 16'b0001100001111110 ; sin_tmp = 16'b0011101100100001 ; end 
  12'd603: begin cos_tmp = 16'b0001100001001110 ; sin_tmp = 16'b0011101100110100 ; end 
  12'd604: begin cos_tmp = 16'b0001100001001110 ; sin_tmp = 16'b0011101100110100 ; end 
  12'd605: begin cos_tmp = 16'b0001100000011111 ; sin_tmp = 16'b0011101101001000 ; end 
  12'd606: begin cos_tmp = 16'b0001011111101111 ; sin_tmp = 16'b0011101101011011 ; end 
  12'd607: begin cos_tmp = 16'b0001011111101111 ; sin_tmp = 16'b0011101101011011 ; end 
  12'd608: begin cos_tmp = 16'b0001011110111111 ; sin_tmp = 16'b0011101101101110 ; end 
  12'd609: begin cos_tmp = 16'b0001011110111111 ; sin_tmp = 16'b0011101101101110 ; end 
  12'd610: begin cos_tmp = 16'b0001011110001111 ; sin_tmp = 16'b0011101110000001 ; end 
  12'd611: begin cos_tmp = 16'b0001011101011111 ; sin_tmp = 16'b0011101110010100 ; end 
  12'd612: begin cos_tmp = 16'b0001011101011111 ; sin_tmp = 16'b0011101110010100 ; end 
  12'd613: begin cos_tmp = 16'b0001011100110000 ; sin_tmp = 16'b0011101110100111 ; end 
  12'd614: begin cos_tmp = 16'b0001011100000000 ; sin_tmp = 16'b0011101110111010 ; end 
  12'd615: begin cos_tmp = 16'b0001011100000000 ; sin_tmp = 16'b0011101110111010 ; end 
  12'd616: begin cos_tmp = 16'b0001011011001111 ; sin_tmp = 16'b0011101111001100 ; end 
  12'd617: begin cos_tmp = 16'b0001011011001111 ; sin_tmp = 16'b0011101111001100 ; end 
  12'd618: begin cos_tmp = 16'b0001011010011111 ; sin_tmp = 16'b0011101111011110 ; end 
  12'd619: begin cos_tmp = 16'b0001011001101111 ; sin_tmp = 16'b0011101111110000 ; end 
  12'd620: begin cos_tmp = 16'b0001011001101111 ; sin_tmp = 16'b0011101111110000 ; end 
  12'd621: begin cos_tmp = 16'b0001011000111111 ; sin_tmp = 16'b0011110000000010 ; end 
  12'd622: begin cos_tmp = 16'b0001011000001111 ; sin_tmp = 16'b0011110000010100 ; end 
  12'd623: begin cos_tmp = 16'b0001011000001111 ; sin_tmp = 16'b0011110000010100 ; end 
  12'd624: begin cos_tmp = 16'b0001010111011110 ; sin_tmp = 16'b0011110000100110 ; end 
  12'd625: begin cos_tmp = 16'b0001010111011110 ; sin_tmp = 16'b0011110000100110 ; end 
  12'd626: begin cos_tmp = 16'b0001010110101110 ; sin_tmp = 16'b0011110000110111 ; end 
  12'd627: begin cos_tmp = 16'b0001010101111101 ; sin_tmp = 16'b0011110001001001 ; end 
  12'd628: begin cos_tmp = 16'b0001010101111101 ; sin_tmp = 16'b0011110001001001 ; end 
  12'd629: begin cos_tmp = 16'b0001010101001101 ; sin_tmp = 16'b0011110001011010 ; end 
  12'd630: begin cos_tmp = 16'b0001010101001101 ; sin_tmp = 16'b0011110001011010 ; end 
  12'd631: begin cos_tmp = 16'b0001010100011100 ; sin_tmp = 16'b0011110001101011 ; end 
  12'd632: begin cos_tmp = 16'b0001010011101100 ; sin_tmp = 16'b0011110001111100 ; end 
  12'd633: begin cos_tmp = 16'b0001010011101100 ; sin_tmp = 16'b0011110001111100 ; end 
  12'd634: begin cos_tmp = 16'b0001010010111011 ; sin_tmp = 16'b0011110010001101 ; end 
  12'd635: begin cos_tmp = 16'b0001010010001010 ; sin_tmp = 16'b0011110010011101 ; end 
  12'd636: begin cos_tmp = 16'b0001010010001010 ; sin_tmp = 16'b0011110010011101 ; end 
  12'd637: begin cos_tmp = 16'b0001010001011010 ; sin_tmp = 16'b0011110010101110 ; end 
  12'd638: begin cos_tmp = 16'b0001010001011010 ; sin_tmp = 16'b0011110010101110 ; end 
  12'd639: begin cos_tmp = 16'b0001010000101001 ; sin_tmp = 16'b0011110010111110 ; end 
  12'd640: begin cos_tmp = 16'b0001001111111000 ; sin_tmp = 16'b0011110011001110 ; end 
  12'd641: begin cos_tmp = 16'b0001001111111000 ; sin_tmp = 16'b0011110011001110 ; end 
  12'd642: begin cos_tmp = 16'b0001001111000111 ; sin_tmp = 16'b0011110011011110 ; end 
  12'd643: begin cos_tmp = 16'b0001001110010110 ; sin_tmp = 16'b0011110011101110 ; end 
  12'd644: begin cos_tmp = 16'b0001001110010110 ; sin_tmp = 16'b0011110011101110 ; end 
  12'd645: begin cos_tmp = 16'b0001001101100101 ; sin_tmp = 16'b0011110011111110 ; end 
  12'd646: begin cos_tmp = 16'b0001001101100101 ; sin_tmp = 16'b0011110011111110 ; end 
  12'd647: begin cos_tmp = 16'b0001001100110100 ; sin_tmp = 16'b0011110100001101 ; end 
  12'd648: begin cos_tmp = 16'b0001001100000011 ; sin_tmp = 16'b0011110100011101 ; end 
  12'd649: begin cos_tmp = 16'b0001001100000011 ; sin_tmp = 16'b0011110100011101 ; end 
  12'd650: begin cos_tmp = 16'b0001001011010010 ; sin_tmp = 16'b0011110100101100 ; end 
  12'd651: begin cos_tmp = 16'b0001001010100000 ; sin_tmp = 16'b0011110100111011 ; end 
  12'd652: begin cos_tmp = 16'b0001001010100000 ; sin_tmp = 16'b0011110100111011 ; end 
  12'd653: begin cos_tmp = 16'b0001001001101111 ; sin_tmp = 16'b0011110101001010 ; end 
  12'd654: begin cos_tmp = 16'b0001001001101111 ; sin_tmp = 16'b0011110101001010 ; end 
  12'd655: begin cos_tmp = 16'b0001001000111110 ; sin_tmp = 16'b0011110101011000 ; end 
  12'd656: begin cos_tmp = 16'b0001001000001100 ; sin_tmp = 16'b0011110101100111 ; end 
  12'd657: begin cos_tmp = 16'b0001001000001100 ; sin_tmp = 16'b0011110101100111 ; end 
  12'd658: begin cos_tmp = 16'b0001000111011011 ; sin_tmp = 16'b0011110101110101 ; end 
  12'd659: begin cos_tmp = 16'b0001000110101010 ; sin_tmp = 16'b0011110110000100 ; end 
  12'd660: begin cos_tmp = 16'b0001000110101010 ; sin_tmp = 16'b0011110110000100 ; end 
  12'd661: begin cos_tmp = 16'b0001000101111000 ; sin_tmp = 16'b0011110110010010 ; end 
  12'd662: begin cos_tmp = 16'b0001000101111000 ; sin_tmp = 16'b0011110110010010 ; end 
  12'd663: begin cos_tmp = 16'b0001000101000111 ; sin_tmp = 16'b0011110110100000 ; end 
  12'd664: begin cos_tmp = 16'b0001000100010101 ; sin_tmp = 16'b0011110110101110 ; end 
  12'd665: begin cos_tmp = 16'b0001000100010101 ; sin_tmp = 16'b0011110110101110 ; end 
  12'd666: begin cos_tmp = 16'b0001000011100011 ; sin_tmp = 16'b0011110110111011 ; end 
  12'd667: begin cos_tmp = 16'b0001000011100011 ; sin_tmp = 16'b0011110110111011 ; end 
  12'd668: begin cos_tmp = 16'b0001000010110010 ; sin_tmp = 16'b0011110111001001 ; end 
  12'd669: begin cos_tmp = 16'b0001000010000000 ; sin_tmp = 16'b0011110111010110 ; end 
  12'd670: begin cos_tmp = 16'b0001000010000000 ; sin_tmp = 16'b0011110111010110 ; end 
  12'd671: begin cos_tmp = 16'b0001000001001110 ; sin_tmp = 16'b0011110111100011 ; end 
  12'd672: begin cos_tmp = 16'b0001000000011100 ; sin_tmp = 16'b0011110111110000 ; end 
  12'd673: begin cos_tmp = 16'b0001000000011100 ; sin_tmp = 16'b0011110111110000 ; end 
  12'd674: begin cos_tmp = 16'b0000111111101011 ; sin_tmp = 16'b0011110111111101 ; end 
  12'd675: begin cos_tmp = 16'b0000111111101011 ; sin_tmp = 16'b0011110111111101 ; end 
  12'd676: begin cos_tmp = 16'b0000111110111001 ; sin_tmp = 16'b0011111000001010 ; end 
  12'd677: begin cos_tmp = 16'b0000111110000111 ; sin_tmp = 16'b0011111000010111 ; end 
  12'd678: begin cos_tmp = 16'b0000111110000111 ; sin_tmp = 16'b0011111000010111 ; end 
  12'd679: begin cos_tmp = 16'b0000111101010101 ; sin_tmp = 16'b0011111000100011 ; end 
  12'd680: begin cos_tmp = 16'b0000111100100011 ; sin_tmp = 16'b0011111000101111 ; end 
  12'd681: begin cos_tmp = 16'b0000111100100011 ; sin_tmp = 16'b0011111000101111 ; end 
  12'd682: begin cos_tmp = 16'b0000111011110001 ; sin_tmp = 16'b0011111000111011 ; end 
  12'd683: begin cos_tmp = 16'b0000111011110001 ; sin_tmp = 16'b0011111000111011 ; end 
  12'd684: begin cos_tmp = 16'b0000111010111111 ; sin_tmp = 16'b0011111001000111 ; end 
  12'd685: begin cos_tmp = 16'b0000111010001101 ; sin_tmp = 16'b0011111001010011 ; end 
  12'd686: begin cos_tmp = 16'b0000111010001101 ; sin_tmp = 16'b0011111001010011 ; end 
  12'd687: begin cos_tmp = 16'b0000111001011010 ; sin_tmp = 16'b0011111001011111 ; end 
  12'd688: begin cos_tmp = 16'b0000111000101000 ; sin_tmp = 16'b0011111001101010 ; end 
  12'd689: begin cos_tmp = 16'b0000111000101000 ; sin_tmp = 16'b0011111001101010 ; end 
  12'd690: begin cos_tmp = 16'b0000110111110110 ; sin_tmp = 16'b0011111001110101 ; end 
  12'd691: begin cos_tmp = 16'b0000110111110110 ; sin_tmp = 16'b0011111001110101 ; end 
  12'd692: begin cos_tmp = 16'b0000110111000100 ; sin_tmp = 16'b0011111010000001 ; end 
  12'd693: begin cos_tmp = 16'b0000110110010010 ; sin_tmp = 16'b0011111010001100 ; end 
  12'd694: begin cos_tmp = 16'b0000110110010010 ; sin_tmp = 16'b0011111010001100 ; end 
  12'd695: begin cos_tmp = 16'b0000110101011111 ; sin_tmp = 16'b0011111010010110 ; end 
  12'd696: begin cos_tmp = 16'b0000110100101101 ; sin_tmp = 16'b0011111010100001 ; end 
  12'd697: begin cos_tmp = 16'b0000110100101101 ; sin_tmp = 16'b0011111010100001 ; end 
  12'd698: begin cos_tmp = 16'b0000110011111010 ; sin_tmp = 16'b0011111010101100 ; end 
  12'd699: begin cos_tmp = 16'b0000110011111010 ; sin_tmp = 16'b0011111010101100 ; end 
  12'd700: begin cos_tmp = 16'b0000110011001000 ; sin_tmp = 16'b0011111010110110 ; end 
  12'd701: begin cos_tmp = 16'b0000110010010110 ; sin_tmp = 16'b0011111011000000 ; end 
  12'd702: begin cos_tmp = 16'b0000110010010110 ; sin_tmp = 16'b0011111011000000 ; end 
  12'd703: begin cos_tmp = 16'b0000110001100011 ; sin_tmp = 16'b0011111011001010 ; end 
  12'd704: begin cos_tmp = 16'b0000110001100011 ; sin_tmp = 16'b0011111011001010 ; end 
  12'd705: begin cos_tmp = 16'b0000110000110001 ; sin_tmp = 16'b0011111011010100 ; end 
  12'd706: begin cos_tmp = 16'b0000101111111110 ; sin_tmp = 16'b0011111011011110 ; end 
  12'd707: begin cos_tmp = 16'b0000101111111110 ; sin_tmp = 16'b0011111011011110 ; end 
  12'd708: begin cos_tmp = 16'b0000101111001011 ; sin_tmp = 16'b0011111011100111 ; end 
  12'd709: begin cos_tmp = 16'b0000101110011001 ; sin_tmp = 16'b0011111011110001 ; end 
  12'd710: begin cos_tmp = 16'b0000101110011001 ; sin_tmp = 16'b0011111011110001 ; end 
  12'd711: begin cos_tmp = 16'b0000101101100110 ; sin_tmp = 16'b0011111011111010 ; end 
  12'd712: begin cos_tmp = 16'b0000101101100110 ; sin_tmp = 16'b0011111011111010 ; end 
  12'd713: begin cos_tmp = 16'b0000101100110100 ; sin_tmp = 16'b0011111100000011 ; end 
  12'd714: begin cos_tmp = 16'b0000101100000001 ; sin_tmp = 16'b0011111100001100 ; end 
  12'd715: begin cos_tmp = 16'b0000101100000001 ; sin_tmp = 16'b0011111100001100 ; end 
  12'd716: begin cos_tmp = 16'b0000101011001110 ; sin_tmp = 16'b0011111100010101 ; end 
  12'd717: begin cos_tmp = 16'b0000101010011011 ; sin_tmp = 16'b0011111100011101 ; end 
  12'd718: begin cos_tmp = 16'b0000101010011011 ; sin_tmp = 16'b0011111100011101 ; end 
  12'd719: begin cos_tmp = 16'b0000101001101001 ; sin_tmp = 16'b0011111100100110 ; end 
  12'd720: begin cos_tmp = 16'b0000101001101001 ; sin_tmp = 16'b0011111100100110 ; end 
  12'd721: begin cos_tmp = 16'b0000101000110110 ; sin_tmp = 16'b0011111100101110 ; end 
  12'd722: begin cos_tmp = 16'b0000101000000011 ; sin_tmp = 16'b0011111100110110 ; end 
  12'd723: begin cos_tmp = 16'b0000101000000011 ; sin_tmp = 16'b0011111100110110 ; end 
  12'd724: begin cos_tmp = 16'b0000100111010000 ; sin_tmp = 16'b0011111100111110 ; end 
  12'd725: begin cos_tmp = 16'b0000100110011101 ; sin_tmp = 16'b0011111101000110 ; end 
  12'd726: begin cos_tmp = 16'b0000100110011101 ; sin_tmp = 16'b0011111101000110 ; end 
  12'd727: begin cos_tmp = 16'b0000100101101010 ; sin_tmp = 16'b0011111101001110 ; end 
  12'd728: begin cos_tmp = 16'b0000100101101010 ; sin_tmp = 16'b0011111101001110 ; end 
  12'd729: begin cos_tmp = 16'b0000100100110111 ; sin_tmp = 16'b0011111101010101 ; end 
  12'd730: begin cos_tmp = 16'b0000100100000101 ; sin_tmp = 16'b0011111101011101 ; end 
  12'd731: begin cos_tmp = 16'b0000100100000101 ; sin_tmp = 16'b0011111101011101 ; end 
  12'd732: begin cos_tmp = 16'b0000100011010010 ; sin_tmp = 16'b0011111101100100 ; end 
  12'd733: begin cos_tmp = 16'b0000100010011111 ; sin_tmp = 16'b0011111101101011 ; end 
  12'd734: begin cos_tmp = 16'b0000100010011111 ; sin_tmp = 16'b0011111101101011 ; end 
  12'd735: begin cos_tmp = 16'b0000100001101100 ; sin_tmp = 16'b0011111101110010 ; end 
  12'd736: begin cos_tmp = 16'b0000100001101100 ; sin_tmp = 16'b0011111101110010 ; end 
  12'd737: begin cos_tmp = 16'b0000100000111001 ; sin_tmp = 16'b0011111101111000 ; end 
  12'd738: begin cos_tmp = 16'b0000100000000101 ; sin_tmp = 16'b0011111101111111 ; end 
  12'd739: begin cos_tmp = 16'b0000100000000101 ; sin_tmp = 16'b0011111101111111 ; end 
  12'd740: begin cos_tmp = 16'b0000011111010010 ; sin_tmp = 16'b0011111110000101 ; end 
  12'd741: begin cos_tmp = 16'b0000011111010010 ; sin_tmp = 16'b0011111110000101 ; end 
  12'd742: begin cos_tmp = 16'b0000011110011111 ; sin_tmp = 16'b0011111110001011 ; end 
  12'd743: begin cos_tmp = 16'b0000011101101100 ; sin_tmp = 16'b0011111110010001 ; end 
  12'd744: begin cos_tmp = 16'b0000011101101100 ; sin_tmp = 16'b0011111110010001 ; end 
  12'd745: begin cos_tmp = 16'b0000011100111001 ; sin_tmp = 16'b0011111110010111 ; end 
  12'd746: begin cos_tmp = 16'b0000011100000110 ; sin_tmp = 16'b0011111110011101 ; end 
  12'd747: begin cos_tmp = 16'b0000011100000110 ; sin_tmp = 16'b0011111110011101 ; end 
  12'd748: begin cos_tmp = 16'b0000011011010011 ; sin_tmp = 16'b0011111110100011 ; end 
  12'd749: begin cos_tmp = 16'b0000011011010011 ; sin_tmp = 16'b0011111110100011 ; end 
  12'd750: begin cos_tmp = 16'b0000011010100000 ; sin_tmp = 16'b0011111110101000 ; end 
  12'd751: begin cos_tmp = 16'b0000011001101100 ; sin_tmp = 16'b0011111110101101 ; end 
  12'd752: begin cos_tmp = 16'b0000011001101100 ; sin_tmp = 16'b0011111110101101 ; end 
  12'd753: begin cos_tmp = 16'b0000011000111001 ; sin_tmp = 16'b0011111110110010 ; end 
  12'd754: begin cos_tmp = 16'b0000011000000110 ; sin_tmp = 16'b0011111110110111 ; end 
  12'd755: begin cos_tmp = 16'b0000011000000110 ; sin_tmp = 16'b0011111110110111 ; end 
  12'd756: begin cos_tmp = 16'b0000010111010011 ; sin_tmp = 16'b0011111110111100 ; end 
  12'd757: begin cos_tmp = 16'b0000010111010011 ; sin_tmp = 16'b0011111110111100 ; end 
  12'd758: begin cos_tmp = 16'b0000010110011111 ; sin_tmp = 16'b0011111111000001 ; end 
  12'd759: begin cos_tmp = 16'b0000010101101100 ; sin_tmp = 16'b0011111111000101 ; end 
  12'd760: begin cos_tmp = 16'b0000010101101100 ; sin_tmp = 16'b0011111111000101 ; end 
  12'd761: begin cos_tmp = 16'b0000010100111001 ; sin_tmp = 16'b0011111111001001 ; end 
  12'd762: begin cos_tmp = 16'b0000010100000101 ; sin_tmp = 16'b0011111111001101 ; end 
  12'd763: begin cos_tmp = 16'b0000010100000101 ; sin_tmp = 16'b0011111111001101 ; end 
  12'd764: begin cos_tmp = 16'b0000010011010010 ; sin_tmp = 16'b0011111111010001 ; end 
  12'd765: begin cos_tmp = 16'b0000010011010010 ; sin_tmp = 16'b0011111111010001 ; end 
  12'd766: begin cos_tmp = 16'b0000010010011111 ; sin_tmp = 16'b0011111111010101 ; end 
  12'd767: begin cos_tmp = 16'b0000010001101011 ; sin_tmp = 16'b0011111111011001 ; end 
  12'd768: begin cos_tmp = 16'b0000010001101011 ; sin_tmp = 16'b0011111111011001 ; end 
  12'd769: begin cos_tmp = 16'b0000010000111000 ; sin_tmp = 16'b0011111111011100 ; end 
  12'd770: begin cos_tmp = 16'b0000010000000101 ; sin_tmp = 16'b0011111111100000 ; end 
  12'd771: begin cos_tmp = 16'b0000010000000101 ; sin_tmp = 16'b0011111111100000 ; end 
  12'd772: begin cos_tmp = 16'b0000001111010001 ; sin_tmp = 16'b0011111111100011 ; end 
  12'd773: begin cos_tmp = 16'b0000001111010001 ; sin_tmp = 16'b0011111111100011 ; end 
  12'd774: begin cos_tmp = 16'b0000001110011110 ; sin_tmp = 16'b0011111111100110 ; end 
  12'd775: begin cos_tmp = 16'b0000001101101011 ; sin_tmp = 16'b0011111111101001 ; end 
  12'd776: begin cos_tmp = 16'b0000001101101011 ; sin_tmp = 16'b0011111111101001 ; end 
  12'd777: begin cos_tmp = 16'b0000001100110111 ; sin_tmp = 16'b0011111111101011 ; end 
  12'd778: begin cos_tmp = 16'b0000001100110111 ; sin_tmp = 16'b0011111111101011 ; end 
  12'd779: begin cos_tmp = 16'b0000001100000100 ; sin_tmp = 16'b0011111111101110 ; end 
  12'd780: begin cos_tmp = 16'b0000001011010000 ; sin_tmp = 16'b0011111111110000 ; end 
  12'd781: begin cos_tmp = 16'b0000001011010000 ; sin_tmp = 16'b0011111111110000 ; end 
  12'd782: begin cos_tmp = 16'b0000001010011101 ; sin_tmp = 16'b0011111111110010 ; end 
  12'd783: begin cos_tmp = 16'b0000001001101010 ; sin_tmp = 16'b0011111111110100 ; end 
  12'd784: begin cos_tmp = 16'b0000001001101010 ; sin_tmp = 16'b0011111111110100 ; end 
  12'd785: begin cos_tmp = 16'b0000001000110110 ; sin_tmp = 16'b0011111111110110 ; end 
  12'd786: begin cos_tmp = 16'b0000001000110110 ; sin_tmp = 16'b0011111111110110 ; end 
  12'd787: begin cos_tmp = 16'b0000001000000011 ; sin_tmp = 16'b0011111111111000 ; end 
  12'd788: begin cos_tmp = 16'b0000000111001111 ; sin_tmp = 16'b0011111111111001 ; end 
  12'd789: begin cos_tmp = 16'b0000000111001111 ; sin_tmp = 16'b0011111111111001 ; end 
  12'd790: begin cos_tmp = 16'b0000000110011100 ; sin_tmp = 16'b0011111111111011 ; end 
  12'd791: begin cos_tmp = 16'b0000000101101000 ; sin_tmp = 16'b0011111111111100 ; end 
  12'd792: begin cos_tmp = 16'b0000000101101000 ; sin_tmp = 16'b0011111111111100 ; end 
  12'd793: begin cos_tmp = 16'b0000000100110101 ; sin_tmp = 16'b0011111111111101 ; end 
  12'd794: begin cos_tmp = 16'b0000000100110101 ; sin_tmp = 16'b0011111111111101 ; end 
  12'd795: begin cos_tmp = 16'b0000000100000001 ; sin_tmp = 16'b0011111111111110 ; end 
  12'd796: begin cos_tmp = 16'b0000000011001110 ; sin_tmp = 16'b0011111111111111 ; end 
  12'd797: begin cos_tmp = 16'b0000000011001110 ; sin_tmp = 16'b0011111111111111 ; end 
  12'd798: begin cos_tmp = 16'b0000000010011010 ; sin_tmp = 16'b0011111111111111 ; end 
  12'd799: begin cos_tmp = 16'b0000000001100111 ; sin_tmp = 16'b0100000000000000 ; end 
  12'd800: begin cos_tmp = 16'b0000000001100111 ; sin_tmp = 16'b0100000000000000 ; end 
  12'd801: begin cos_tmp = 16'b0000000000110011 ; sin_tmp = 16'b0100000000000000 ; end 
  12'd802: begin cos_tmp = 16'b0000000000110011 ; sin_tmp = 16'b0100000000000000 ; end 
  12'd803: begin cos_tmp = 16'b0000000000000000 ; sin_tmp = 16'b0100000000000000 ; end 
  endcase
end
endmodule
